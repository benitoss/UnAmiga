-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80e4",
     9 => x"b4080b0b",
    10 => x"80e4b808",
    11 => x"0b0b80e4",
    12 => x"bc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"e4bc0c0b",
    16 => x"0b80e4b8",
    17 => x"0c0b0b80",
    18 => x"e4b40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80dfa4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80e4b470",
    57 => x"80eef027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51b192",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80e4",
    65 => x"c40c9f0b",
    66 => x"80e4c80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"e4c808ff",
    70 => x"0580e4c8",
    71 => x"0c80e4c8",
    72 => x"088025e8",
    73 => x"3880e4c4",
    74 => x"08ff0580",
    75 => x"e4c40c80",
    76 => x"e4c40880",
    77 => x"25d03880",
    78 => x"0b80e4c8",
    79 => x"0c800b80",
    80 => x"e4c40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80e4c408",
   100 => x"25913882",
   101 => x"c82d80e4",
   102 => x"c408ff05",
   103 => x"80e4c40c",
   104 => x"838a0480",
   105 => x"e4c40880",
   106 => x"e4c80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80e4c408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"e4c80881",
   116 => x"0580e4c8",
   117 => x"0c80e4c8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80e4c8",
   121 => x"0c80e4c4",
   122 => x"08810580",
   123 => x"e4c40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480e4",
   128 => x"c8088105",
   129 => x"80e4c80c",
   130 => x"80e4c808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80e4c8",
   134 => x"0c80e4c4",
   135 => x"08810580",
   136 => x"e4c40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"e4cc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"e4cc0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280e4",
   177 => x"cc088407",
   178 => x"80e4cc0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80e1",
   183 => x"c40c8171",
   184 => x"2bff05f6",
   185 => x"880cfdfc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80e4cc",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80e4",
   208 => x"b40c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"a00bec0c",
  1093 => x"86c72d86",
  1094 => x"c72d86c7",
  1095 => x"2d86c72d",
  1096 => x"86c72d86",
  1097 => x"c72d86c7",
  1098 => x"2d86c72d",
  1099 => x"86c72d86",
  1100 => x"c72d86c7",
  1101 => x"2d86c72d",
  1102 => x"86c72d86",
  1103 => x"c72d86c7",
  1104 => x"2d86c72d",
  1105 => x"86c72d86",
  1106 => x"c72d86c7",
  1107 => x"2d86c72d",
  1108 => x"86c72d86",
  1109 => x"c72d86c7",
  1110 => x"2d86c72d",
  1111 => x"86c72d86",
  1112 => x"c72d86c7",
  1113 => x"2d86c72d",
  1114 => x"86c72d86",
  1115 => x"c72d86c7",
  1116 => x"2d86c72d",
  1117 => x"86c72d86",
  1118 => x"c72d86c7",
  1119 => x"2d86c72d",
  1120 => x"86c72d86",
  1121 => x"c72d86c7",
  1122 => x"2d86c72d",
  1123 => x"86c72d86",
  1124 => x"c72d86c7",
  1125 => x"2d86c72d",
  1126 => x"86c72d86",
  1127 => x"c72d86c7",
  1128 => x"2d86c72d",
  1129 => x"86c72d86",
  1130 => x"c72d86c7",
  1131 => x"2d86c72d",
  1132 => x"86c72d86",
  1133 => x"c72d86c7",
  1134 => x"2d86c72d",
  1135 => x"86c72d86",
  1136 => x"c72d86c7",
  1137 => x"2d86c72d",
  1138 => x"86c72d86",
  1139 => x"c72d86c7",
  1140 => x"2d86c72d",
  1141 => x"86c72d86",
  1142 => x"c72d86c7",
  1143 => x"2d86c72d",
  1144 => x"86c72d86",
  1145 => x"c72d86c7",
  1146 => x"2d86c72d",
  1147 => x"86c72d86",
  1148 => x"c72d86c7",
  1149 => x"2d86c72d",
  1150 => x"86c72d86",
  1151 => x"c72d86c7",
  1152 => x"2d86c72d",
  1153 => x"86c72d86",
  1154 => x"c72d86c7",
  1155 => x"2d86c72d",
  1156 => x"86c72d86",
  1157 => x"c72d86c7",
  1158 => x"2d86c72d",
  1159 => x"86c72d86",
  1160 => x"c72d86c7",
  1161 => x"2d86c72d",
  1162 => x"86c72d86",
  1163 => x"c72d86c7",
  1164 => x"2d86c72d",
  1165 => x"86c72d86",
  1166 => x"c72d86c7",
  1167 => x"2d86c72d",
  1168 => x"86c72d86",
  1169 => x"c72d86c7",
  1170 => x"2d86c72d",
  1171 => x"86c72d86",
  1172 => x"c72d86c7",
  1173 => x"2d86c72d",
  1174 => x"86c72d86",
  1175 => x"c72d86c7",
  1176 => x"2d86c72d",
  1177 => x"86c72d86",
  1178 => x"c72d86c7",
  1179 => x"2d86c72d",
  1180 => x"86c72d86",
  1181 => x"c72d86c7",
  1182 => x"2d86c72d",
  1183 => x"86c72d86",
  1184 => x"c72d86c7",
  1185 => x"2d86c72d",
  1186 => x"86c72d86",
  1187 => x"c72d86c7",
  1188 => x"2d86c72d",
  1189 => x"86c72d86",
  1190 => x"c72d86c7",
  1191 => x"2d86c72d",
  1192 => x"86c72d86",
  1193 => x"c72d86c7",
  1194 => x"2d86c72d",
  1195 => x"86c72d86",
  1196 => x"c72d86c7",
  1197 => x"2d86c72d",
  1198 => x"86c72d86",
  1199 => x"c72d86c7",
  1200 => x"2d86c72d",
  1201 => x"86c72d86",
  1202 => x"c72d86c7",
  1203 => x"2d86c72d",
  1204 => x"86c72d86",
  1205 => x"c72d86c7",
  1206 => x"2d86c72d",
  1207 => x"86c72d86",
  1208 => x"c72d86c7",
  1209 => x"2d86c72d",
  1210 => x"86c72d86",
  1211 => x"c72d86c7",
  1212 => x"2d86c72d",
  1213 => x"86c72d86",
  1214 => x"c72d86c7",
  1215 => x"2d86c72d",
  1216 => x"86c72d86",
  1217 => x"c72d86c7",
  1218 => x"2d86c72d",
  1219 => x"86c72d86",
  1220 => x"c72d86c7",
  1221 => x"2d86c72d",
  1222 => x"86c72d86",
  1223 => x"c72d86c7",
  1224 => x"2d86c72d",
  1225 => x"86c72d86",
  1226 => x"c72d86c7",
  1227 => x"2d86c72d",
  1228 => x"86c72d86",
  1229 => x"c72d86c7",
  1230 => x"2d86c72d",
  1231 => x"86c72d86",
  1232 => x"c72d86c7",
  1233 => x"2d86c72d",
  1234 => x"86c72d86",
  1235 => x"c72d86c7",
  1236 => x"2d86c72d",
  1237 => x"86c72d86",
  1238 => x"c72d86c7",
  1239 => x"2d86c72d",
  1240 => x"86c72d86",
  1241 => x"c72d86c7",
  1242 => x"2d86c72d",
  1243 => x"86c72d86",
  1244 => x"c72d86c7",
  1245 => x"2d86c72d",
  1246 => x"86c72d86",
  1247 => x"c72d86c7",
  1248 => x"2d86c72d",
  1249 => x"86c72d86",
  1250 => x"c72d86c7",
  1251 => x"2d86c72d",
  1252 => x"86c72d86",
  1253 => x"c72d86c7",
  1254 => x"2d86c72d",
  1255 => x"86c72d86",
  1256 => x"c72d86c7",
  1257 => x"2d86c72d",
  1258 => x"86c72d86",
  1259 => x"c72d86c7",
  1260 => x"2d86c72d",
  1261 => x"86c72d86",
  1262 => x"c72d86c7",
  1263 => x"2d86c72d",
  1264 => x"86c72d86",
  1265 => x"c72d86c7",
  1266 => x"2d86c72d",
  1267 => x"86c72d86",
  1268 => x"c72d86c7",
  1269 => x"2d86c72d",
  1270 => x"86c72d86",
  1271 => x"c72d86c7",
  1272 => x"2d86c72d",
  1273 => x"86c72d86",
  1274 => x"c72d86c7",
  1275 => x"2d86c72d",
  1276 => x"86c72d86",
  1277 => x"c72d86c7",
  1278 => x"2d86c72d",
  1279 => x"86c72d86",
  1280 => x"c72d86c7",
  1281 => x"2d86c72d",
  1282 => x"86c72d86",
  1283 => x"c72d86c7",
  1284 => x"2d86c72d",
  1285 => x"86c72d86",
  1286 => x"c72d86c7",
  1287 => x"2d86c72d",
  1288 => x"86c72d86",
  1289 => x"c72d86c7",
  1290 => x"2d86c72d",
  1291 => x"86c72d86",
  1292 => x"c72d86c7",
  1293 => x"2d86c72d",
  1294 => x"86c72d86",
  1295 => x"c72d86c7",
  1296 => x"2d86c72d",
  1297 => x"86c72d86",
  1298 => x"c72d86c7",
  1299 => x"2d86c72d",
  1300 => x"86c72d86",
  1301 => x"c72d86c7",
  1302 => x"2d86c72d",
  1303 => x"86c72d86",
  1304 => x"c72d86c7",
  1305 => x"2d86c72d",
  1306 => x"86c72d86",
  1307 => x"c72d86c7",
  1308 => x"2d86c72d",
  1309 => x"86c72d86",
  1310 => x"c72d86c7",
  1311 => x"2d86c72d",
  1312 => x"86c72d86",
  1313 => x"c72d86c7",
  1314 => x"2d86c72d",
  1315 => x"86c72d86",
  1316 => x"c72d86c7",
  1317 => x"2d86c72d",
  1318 => x"86c72d86",
  1319 => x"c72d86c7",
  1320 => x"2d86c72d",
  1321 => x"86c72d86",
  1322 => x"c72d86c7",
  1323 => x"2d86c72d",
  1324 => x"86c72d86",
  1325 => x"c72d86c7",
  1326 => x"2d86c72d",
  1327 => x"86c72d86",
  1328 => x"c72d86c7",
  1329 => x"2d86c72d",
  1330 => x"86c72d86",
  1331 => x"c72d86c7",
  1332 => x"2d86c72d",
  1333 => x"86c72d86",
  1334 => x"c72d86c7",
  1335 => x"2d86c72d",
  1336 => x"86c72d86",
  1337 => x"c72d86c7",
  1338 => x"2d86c72d",
  1339 => x"86c72d86",
  1340 => x"c72d86c7",
  1341 => x"2d86c72d",
  1342 => x"86c72d86",
  1343 => x"c72d86c7",
  1344 => x"2d86c72d",
  1345 => x"86c72d86",
  1346 => x"c72d86c7",
  1347 => x"2d86c72d",
  1348 => x"86c72d86",
  1349 => x"c72d86c7",
  1350 => x"2d86c72d",
  1351 => x"86c72d86",
  1352 => x"c72d86c7",
  1353 => x"2d86c72d",
  1354 => x"86c72d86",
  1355 => x"c72d86c7",
  1356 => x"2d86c72d",
  1357 => x"86c72d86",
  1358 => x"c72d86c7",
  1359 => x"2d86c72d",
  1360 => x"86c72d86",
  1361 => x"c72d86c7",
  1362 => x"2d86c72d",
  1363 => x"86c72d86",
  1364 => x"c72d86c7",
  1365 => x"2d86c72d",
  1366 => x"86c72d86",
  1367 => x"c72d86c7",
  1368 => x"2d86c72d",
  1369 => x"86c72d86",
  1370 => x"c72d86c7",
  1371 => x"2d86c72d",
  1372 => x"86c72d86",
  1373 => x"c72d86c7",
  1374 => x"2d86c72d",
  1375 => x"86c72d86",
  1376 => x"c72d86c7",
  1377 => x"2d86c72d",
  1378 => x"86c72d86",
  1379 => x"c72d86c7",
  1380 => x"2d86c72d",
  1381 => x"86c72d86",
  1382 => x"c72d86c7",
  1383 => x"2d86c72d",
  1384 => x"86c72d86",
  1385 => x"c72d86c7",
  1386 => x"2d86c72d",
  1387 => x"86c72d86",
  1388 => x"c72d86c7",
  1389 => x"2d86c72d",
  1390 => x"86c72d86",
  1391 => x"c72d86c7",
  1392 => x"2d86c72d",
  1393 => x"86c72d86",
  1394 => x"c72d86c7",
  1395 => x"2d86c72d",
  1396 => x"86c72d86",
  1397 => x"c72d86c7",
  1398 => x"2d86c72d",
  1399 => x"86c72d86",
  1400 => x"c72d86c7",
  1401 => x"2d86c72d",
  1402 => x"86c72d86",
  1403 => x"c72d86c7",
  1404 => x"2d86c72d",
  1405 => x"86c72d86",
  1406 => x"c72d86c7",
  1407 => x"2d86c72d",
  1408 => x"86c72d86",
  1409 => x"c72d86c7",
  1410 => x"2d86c72d",
  1411 => x"86c72d86",
  1412 => x"c72d86c7",
  1413 => x"2d86c72d",
  1414 => x"86c72d86",
  1415 => x"c72d86c7",
  1416 => x"2d86c72d",
  1417 => x"86c72d86",
  1418 => x"c72d86c7",
  1419 => x"2d86c72d",
  1420 => x"86c72d86",
  1421 => x"c72d86c7",
  1422 => x"2d86c72d",
  1423 => x"86c72d86",
  1424 => x"c72d86c7",
  1425 => x"2d86c72d",
  1426 => x"86c72d86",
  1427 => x"c72d86c7",
  1428 => x"2d86c72d",
  1429 => x"86c72d86",
  1430 => x"c72d86c7",
  1431 => x"2d86c72d",
  1432 => x"86c72d86",
  1433 => x"c72d86c7",
  1434 => x"2d86c72d",
  1435 => x"86c72d86",
  1436 => x"c72d86c7",
  1437 => x"2d86c72d",
  1438 => x"86c72d86",
  1439 => x"c72d86c7",
  1440 => x"2d86c72d",
  1441 => x"86c72d86",
  1442 => x"c72d86c7",
  1443 => x"2d86c72d",
  1444 => x"86c72d86",
  1445 => x"c72d86c7",
  1446 => x"2d86c72d",
  1447 => x"86c72d86",
  1448 => x"c72d86c7",
  1449 => x"2d86c72d",
  1450 => x"86c72d86",
  1451 => x"c72d86c7",
  1452 => x"2d86c72d",
  1453 => x"86c72d86",
  1454 => x"c72d86c7",
  1455 => x"2d86c72d",
  1456 => x"86c72d86",
  1457 => x"c72d86c7",
  1458 => x"2d86c72d",
  1459 => x"86c72d86",
  1460 => x"c72d86c7",
  1461 => x"2d86c72d",
  1462 => x"86c72d86",
  1463 => x"c72d86c7",
  1464 => x"2d86c72d",
  1465 => x"86c72d86",
  1466 => x"c72d86c7",
  1467 => x"2d86c72d",
  1468 => x"86c72d86",
  1469 => x"c72d86c7",
  1470 => x"2d86c72d",
  1471 => x"86c72d86",
  1472 => x"c72d86c7",
  1473 => x"2d86c72d",
  1474 => x"86c72d86",
  1475 => x"c72d86c7",
  1476 => x"2d86c72d",
  1477 => x"86c72d86",
  1478 => x"c72d86c7",
  1479 => x"2d86c72d",
  1480 => x"86c72d86",
  1481 => x"c72d86c7",
  1482 => x"2d86c72d",
  1483 => x"86c72d86",
  1484 => x"c72d86c7",
  1485 => x"2d86c72d",
  1486 => x"86c72d86",
  1487 => x"c72d86c7",
  1488 => x"2d86c72d",
  1489 => x"86c72d86",
  1490 => x"c72d86c7",
  1491 => x"2d86c72d",
  1492 => x"86c72d86",
  1493 => x"c72d86c7",
  1494 => x"2d86c72d",
  1495 => x"86c72d86",
  1496 => x"c72d86c7",
  1497 => x"2d86c72d",
  1498 => x"86c72d86",
  1499 => x"c72d86c7",
  1500 => x"2d86c72d",
  1501 => x"86c72d86",
  1502 => x"c72d86c7",
  1503 => x"2d86c72d",
  1504 => x"86c72d86",
  1505 => x"c72d86c7",
  1506 => x"2d86c72d",
  1507 => x"86c72d86",
  1508 => x"c72d86c7",
  1509 => x"2d86c72d",
  1510 => x"86c72d86",
  1511 => x"c72d86c7",
  1512 => x"2d86c72d",
  1513 => x"86c72d86",
  1514 => x"c72d86c7",
  1515 => x"2d86c72d",
  1516 => x"86c72d86",
  1517 => x"c72d86c7",
  1518 => x"2d86c72d",
  1519 => x"86c72d86",
  1520 => x"c72d86c7",
  1521 => x"2d86c72d",
  1522 => x"86c72d86",
  1523 => x"c72d86c7",
  1524 => x"2d86c72d",
  1525 => x"0402dc05",
  1526 => x"0d8059a2",
  1527 => x"902d810b",
  1528 => x"ec0c7a52",
  1529 => x"80e4d051",
  1530 => x"80d5ef2d",
  1531 => x"80e4b408",
  1532 => x"792e80f7",
  1533 => x"3880e4d4",
  1534 => x"0870f80c",
  1535 => x"79ff1256",
  1536 => x"59557379",
  1537 => x"2e8b3881",
  1538 => x"1874812a",
  1539 => x"555873f7",
  1540 => x"38f71858",
  1541 => x"81598075",
  1542 => x"2580d038",
  1543 => x"77527351",
  1544 => x"84a82d80",
  1545 => x"e5a85280",
  1546 => x"e4d05180",
  1547 => x"d8c52d80",
  1548 => x"e4b40880",
  1549 => x"2e9b3880",
  1550 => x"e5a85783",
  1551 => x"fc567670",
  1552 => x"84055808",
  1553 => x"e80cfc16",
  1554 => x"56758025",
  1555 => x"f138b0d9",
  1556 => x"0480e4b4",
  1557 => x"08598480",
  1558 => x"5580e4d0",
  1559 => x"5180d894",
  1560 => x"2dfc8015",
  1561 => x"81155555",
  1562 => x"b0960484",
  1563 => x"0bec0c78",
  1564 => x"802e8e38",
  1565 => x"80e1c851",
  1566 => x"b8e52db6",
  1567 => x"d82db188",
  1568 => x"0480e284",
  1569 => x"51b8e52d",
  1570 => x"7880e4b4",
  1571 => x"0c02a405",
  1572 => x"0d0402f0",
  1573 => x"050d840b",
  1574 => x"ec0cb68b",
  1575 => x"2db2b92d",
  1576 => x"81f92d83",
  1577 => x"52b5ee2d",
  1578 => x"8151858d",
  1579 => x"2dff1252",
  1580 => x"718025f1",
  1581 => x"38840bec",
  1582 => x"0c80dff8",
  1583 => x"5186a02d",
  1584 => x"80cc8f2d",
  1585 => x"80e4b408",
  1586 => x"802e80d6",
  1587 => x"38afd551",
  1588 => x"80df9c2d",
  1589 => x"80e1c851",
  1590 => x"b8e52db6",
  1591 => x"c42db2c5",
  1592 => x"2db8f82d",
  1593 => x"80e1dc0b",
  1594 => x"80f52d80",
  1595 => x"e2f00870",
  1596 => x"81065455",
  1597 => x"5371802e",
  1598 => x"85387281",
  1599 => x"07537381",
  1600 => x"2a708106",
  1601 => x"51527180",
  1602 => x"2e853872",
  1603 => x"82075372",
  1604 => x"fc0c8652",
  1605 => x"80e4b408",
  1606 => x"83388452",
  1607 => x"71ec0cb1",
  1608 => x"de04800b",
  1609 => x"80e4b40c",
  1610 => x"0290050d",
  1611 => x"0471980c",
  1612 => x"04ffb008",
  1613 => x"80e4b40c",
  1614 => x"04810bff",
  1615 => x"b00c0480",
  1616 => x"0bffb00c",
  1617 => x"0402f405",
  1618 => x"0d80e4dc",
  1619 => x"51b4d82d",
  1620 => x"ff0b80e4",
  1621 => x"b4082581",
  1622 => x"883880e4",
  1623 => x"b40881f0",
  1624 => x"2e098106",
  1625 => x"8a38810b",
  1626 => x"80e2e80c",
  1627 => x"b3e10480",
  1628 => x"e4b40881",
  1629 => x"e02e0981",
  1630 => x"068a3881",
  1631 => x"0b80e2ec",
  1632 => x"0cb3e104",
  1633 => x"80e4b408",
  1634 => x"5280e2ec",
  1635 => x"08802e89",
  1636 => x"3880e4b4",
  1637 => x"08818005",
  1638 => x"5271842c",
  1639 => x"728f0653",
  1640 => x"5380e2e8",
  1641 => x"08802e9a",
  1642 => x"38728429",
  1643 => x"80e2a805",
  1644 => x"72138171",
  1645 => x"2b700973",
  1646 => x"0806730c",
  1647 => x"515353b3",
  1648 => x"d5047284",
  1649 => x"2980e2a8",
  1650 => x"05721383",
  1651 => x"712b7208",
  1652 => x"07720c53",
  1653 => x"53800b80",
  1654 => x"e2ec0c80",
  1655 => x"0b80e2e8",
  1656 => x"0c800b80",
  1657 => x"e4b40c02",
  1658 => x"8c050d04",
  1659 => x"02f8050d",
  1660 => x"80e2a852",
  1661 => x"8f518072",
  1662 => x"70840554",
  1663 => x"0cff1151",
  1664 => x"708025f2",
  1665 => x"38028805",
  1666 => x"0d0402f0",
  1667 => x"050d7551",
  1668 => x"b2bf2d70",
  1669 => x"822cfc06",
  1670 => x"80e2a811",
  1671 => x"72109e06",
  1672 => x"71087072",
  1673 => x"2a708306",
  1674 => x"82742b70",
  1675 => x"09740676",
  1676 => x"0c545156",
  1677 => x"57535153",
  1678 => x"b2b92d71",
  1679 => x"80e4b40c",
  1680 => x"0290050d",
  1681 => x"0402fc05",
  1682 => x"0d725180",
  1683 => x"710c800b",
  1684 => x"84120c02",
  1685 => x"84050d04",
  1686 => x"02f0050d",
  1687 => x"75700884",
  1688 => x"12085353",
  1689 => x"53ff5471",
  1690 => x"712ea838",
  1691 => x"b2bf2d84",
  1692 => x"13087084",
  1693 => x"29148811",
  1694 => x"70087081",
  1695 => x"ff068418",
  1696 => x"08811187",
  1697 => x"06841a0c",
  1698 => x"53515551",
  1699 => x"5151b2b9",
  1700 => x"2d715473",
  1701 => x"80e4b40c",
  1702 => x"0290050d",
  1703 => x"0402f405",
  1704 => x"0db2bf2d",
  1705 => x"e008708b",
  1706 => x"2a708106",
  1707 => x"51525370",
  1708 => x"802ea138",
  1709 => x"80e4dc08",
  1710 => x"70842980",
  1711 => x"e4e40574",
  1712 => x"81ff0671",
  1713 => x"0c515180",
  1714 => x"e4dc0881",
  1715 => x"11870680",
  1716 => x"e4dc0c51",
  1717 => x"728c2cbf",
  1718 => x"0680e584",
  1719 => x"0c800b80",
  1720 => x"e5880cb2",
  1721 => x"b12db2b9",
  1722 => x"2d028c05",
  1723 => x"0d0402fc",
  1724 => x"050db2bf",
  1725 => x"2d810b80",
  1726 => x"e5880cb2",
  1727 => x"b92d80e5",
  1728 => x"88085170",
  1729 => x"f9380284",
  1730 => x"050d0402",
  1731 => x"fc050d80",
  1732 => x"e4dc51b4",
  1733 => x"c52db3ec",
  1734 => x"2db59d51",
  1735 => x"b2ad2d02",
  1736 => x"84050d04",
  1737 => x"02fc050d",
  1738 => x"8fcf5186",
  1739 => x"c72dff11",
  1740 => x"51708025",
  1741 => x"f6380284",
  1742 => x"050d0480",
  1743 => x"e5940880",
  1744 => x"e4b40c04",
  1745 => x"02fc050d",
  1746 => x"810b80e2",
  1747 => x"f40c8151",
  1748 => x"858d2d02",
  1749 => x"84050d04",
  1750 => x"02fc050d",
  1751 => x"b6e204b2",
  1752 => x"c52d80f6",
  1753 => x"51b48a2d",
  1754 => x"80e4b408",
  1755 => x"f23880da",
  1756 => x"51b48a2d",
  1757 => x"80e4b408",
  1758 => x"e63880e4",
  1759 => x"b40880e2",
  1760 => x"f40c80e4",
  1761 => x"b4085185",
  1762 => x"8d2d0284",
  1763 => x"050d0402",
  1764 => x"ec050d76",
  1765 => x"54805287",
  1766 => x"0b881580",
  1767 => x"f52d5653",
  1768 => x"74722483",
  1769 => x"38a05372",
  1770 => x"5183842d",
  1771 => x"81128b15",
  1772 => x"80f52d54",
  1773 => x"52727225",
  1774 => x"de380294",
  1775 => x"050d0402",
  1776 => x"f0050d80",
  1777 => x"e5940854",
  1778 => x"81f92d80",
  1779 => x"0b80e598",
  1780 => x"0c730880",
  1781 => x"2e818938",
  1782 => x"820b80e4",
  1783 => x"c80c80e5",
  1784 => x"98088f06",
  1785 => x"80e4c40c",
  1786 => x"73085271",
  1787 => x"832e9638",
  1788 => x"71832689",
  1789 => x"3871812e",
  1790 => x"b038b8c9",
  1791 => x"0471852e",
  1792 => x"a038b8c9",
  1793 => x"04881480",
  1794 => x"f52d8415",
  1795 => x"0880e090",
  1796 => x"53545286",
  1797 => x"a02d7184",
  1798 => x"29137008",
  1799 => x"5252b8cd",
  1800 => x"047351b7",
  1801 => x"8f2db8c9",
  1802 => x"0480e2f0",
  1803 => x"08881508",
  1804 => x"2c708106",
  1805 => x"51527180",
  1806 => x"2e883880",
  1807 => x"e09451b8",
  1808 => x"c60480e0",
  1809 => x"985186a0",
  1810 => x"2d841408",
  1811 => x"5186a02d",
  1812 => x"80e59808",
  1813 => x"810580e5",
  1814 => x"980c8c14",
  1815 => x"54b7d104",
  1816 => x"0290050d",
  1817 => x"047180e5",
  1818 => x"940cb7bf",
  1819 => x"2d80e598",
  1820 => x"08ff0580",
  1821 => x"e59c0c04",
  1822 => x"02e8050d",
  1823 => x"80e59408",
  1824 => x"80e5a008",
  1825 => x"575580f6",
  1826 => x"51b48a2d",
  1827 => x"80e4b408",
  1828 => x"812a7081",
  1829 => x"06515271",
  1830 => x"802ea238",
  1831 => x"b9a204b2",
  1832 => x"c52d80f6",
  1833 => x"51b48a2d",
  1834 => x"80e4b408",
  1835 => x"f23880e2",
  1836 => x"f4088132",
  1837 => x"7080e2f4",
  1838 => x"0c51858d",
  1839 => x"2d80e584",
  1840 => x"08a00652",
  1841 => x"80722598",
  1842 => x"38b6a42d",
  1843 => x"b2c52d80",
  1844 => x"e2f40881",
  1845 => x"327080e2",
  1846 => x"f40c7052",
  1847 => x"52858d2d",
  1848 => x"800b80e5",
  1849 => x"8c0c800b",
  1850 => x"80e5900c",
  1851 => x"80e2f408",
  1852 => x"83ae3880",
  1853 => x"da51b48a",
  1854 => x"2d80e4b4",
  1855 => x"08802e8c",
  1856 => x"3880e58c",
  1857 => x"08818007",
  1858 => x"80e58c0c",
  1859 => x"80d951b4",
  1860 => x"8a2d80e4",
  1861 => x"b408802e",
  1862 => x"8c3880e5",
  1863 => x"8c0880c0",
  1864 => x"0780e58c",
  1865 => x"0c819451",
  1866 => x"b48a2d80",
  1867 => x"e4b40880",
  1868 => x"2e8b3880",
  1869 => x"e58c0890",
  1870 => x"0780e58c",
  1871 => x"0c819151",
  1872 => x"b48a2d80",
  1873 => x"e4b40880",
  1874 => x"2e8b3880",
  1875 => x"e58c08a0",
  1876 => x"0780e58c",
  1877 => x"0c81f551",
  1878 => x"b48a2d80",
  1879 => x"e4b40880",
  1880 => x"2e8b3880",
  1881 => x"e58c0881",
  1882 => x"0780e58c",
  1883 => x"0c81f251",
  1884 => x"b48a2d80",
  1885 => x"e4b40880",
  1886 => x"2e8b3880",
  1887 => x"e58c0882",
  1888 => x"0780e58c",
  1889 => x"0c81eb51",
  1890 => x"b48a2d80",
  1891 => x"e4b40880",
  1892 => x"2e8b3880",
  1893 => x"e58c0884",
  1894 => x"0780e58c",
  1895 => x"0c81f451",
  1896 => x"b48a2d80",
  1897 => x"e4b40880",
  1898 => x"2e8b3880",
  1899 => x"e58c0888",
  1900 => x"0780e58c",
  1901 => x"0c80d851",
  1902 => x"b48a2d80",
  1903 => x"e4b40880",
  1904 => x"2e8c3880",
  1905 => x"e5900881",
  1906 => x"800780e5",
  1907 => x"900c9251",
  1908 => x"b48a2d80",
  1909 => x"e4b40880",
  1910 => x"2e8c3880",
  1911 => x"e5900880",
  1912 => x"c00780e5",
  1913 => x"900c9451",
  1914 => x"b48a2d80",
  1915 => x"e4b40880",
  1916 => x"2e8b3880",
  1917 => x"e5900890",
  1918 => x"0780e590",
  1919 => x"0c9151b4",
  1920 => x"8a2d80e4",
  1921 => x"b408802e",
  1922 => x"8b3880e5",
  1923 => x"9008a007",
  1924 => x"80e5900c",
  1925 => x"9d51b48a",
  1926 => x"2d80e4b4",
  1927 => x"08802e8b",
  1928 => x"3880e590",
  1929 => x"08810780",
  1930 => x"e5900c9b",
  1931 => x"51b48a2d",
  1932 => x"80e4b408",
  1933 => x"802e8b38",
  1934 => x"80e59008",
  1935 => x"820780e5",
  1936 => x"900c9c51",
  1937 => x"b48a2d80",
  1938 => x"e4b40880",
  1939 => x"2e8b3880",
  1940 => x"e5900884",
  1941 => x"0780e590",
  1942 => x"0ca351b4",
  1943 => x"8a2d80e4",
  1944 => x"b408802e",
  1945 => x"8b3880e5",
  1946 => x"90088807",
  1947 => x"80e5900c",
  1948 => x"9651b48a",
  1949 => x"2d80e4b4",
  1950 => x"08802e84",
  1951 => x"3894bf2d",
  1952 => x"9e51b48a",
  1953 => x"2d80e4b4",
  1954 => x"08802e84",
  1955 => x"3886ee2d",
  1956 => x"81fd51b4",
  1957 => x"8a2d81fa",
  1958 => x"51b48a2d",
  1959 => x"80c3c804",
  1960 => x"81f551b4",
  1961 => x"8a2d80e4",
  1962 => x"b408812a",
  1963 => x"70810651",
  1964 => x"52718e38",
  1965 => x"80e58408",
  1966 => x"90065280",
  1967 => x"722580c2",
  1968 => x"3880e584",
  1969 => x"08900652",
  1970 => x"80722584",
  1971 => x"38b6a42d",
  1972 => x"80e59c08",
  1973 => x"5271802e",
  1974 => x"8a38ff12",
  1975 => x"80e59c0c",
  1976 => x"be820480",
  1977 => x"e5980810",
  1978 => x"80e59808",
  1979 => x"05708429",
  1980 => x"16515288",
  1981 => x"1208802e",
  1982 => x"8938ff51",
  1983 => x"88120852",
  1984 => x"712d81f2",
  1985 => x"51b48a2d",
  1986 => x"80e4b408",
  1987 => x"812a7081",
  1988 => x"06515271",
  1989 => x"8e3880e5",
  1990 => x"84088806",
  1991 => x"52807225",
  1992 => x"80c33880",
  1993 => x"e5840888",
  1994 => x"06528072",
  1995 => x"258438b6",
  1996 => x"a42d80e5",
  1997 => x"9808ff11",
  1998 => x"80e59c08",
  1999 => x"56535373",
  2000 => x"72258a38",
  2001 => x"811480e5",
  2002 => x"9c0cbee5",
  2003 => x"04721013",
  2004 => x"70842916",
  2005 => x"51528812",
  2006 => x"08802e89",
  2007 => x"38fe5188",
  2008 => x"12085271",
  2009 => x"2d81fd51",
  2010 => x"b48a2d80",
  2011 => x"e4b40881",
  2012 => x"2a708106",
  2013 => x"51527180",
  2014 => x"2eb13880",
  2015 => x"e59c0880",
  2016 => x"2e8a3880",
  2017 => x"0b80e59c",
  2018 => x"0cbfab04",
  2019 => x"80e59808",
  2020 => x"1080e598",
  2021 => x"08057084",
  2022 => x"29165152",
  2023 => x"88120880",
  2024 => x"2e8938fd",
  2025 => x"51881208",
  2026 => x"52712d81",
  2027 => x"fa51b48a",
  2028 => x"2d80e4b4",
  2029 => x"08812a70",
  2030 => x"81065152",
  2031 => x"71802eb1",
  2032 => x"3880e598",
  2033 => x"08ff1154",
  2034 => x"5280e59c",
  2035 => x"08732589",
  2036 => x"387280e5",
  2037 => x"9c0cbff1",
  2038 => x"04711012",
  2039 => x"70842916",
  2040 => x"51528812",
  2041 => x"08802e89",
  2042 => x"38fc5188",
  2043 => x"12085271",
  2044 => x"2d80e59c",
  2045 => x"08705354",
  2046 => x"73802e8a",
  2047 => x"388c15ff",
  2048 => x"155555bf",
  2049 => x"f804820b",
  2050 => x"80e4c80c",
  2051 => x"718f0680",
  2052 => x"e4c40c81",
  2053 => x"eb51b48a",
  2054 => x"2d80e4b4",
  2055 => x"08812a70",
  2056 => x"81065152",
  2057 => x"71802ead",
  2058 => x"38740885",
  2059 => x"2e098106",
  2060 => x"a4388815",
  2061 => x"80f52dff",
  2062 => x"05527188",
  2063 => x"1681b72d",
  2064 => x"71982b52",
  2065 => x"71802588",
  2066 => x"38800b88",
  2067 => x"1681b72d",
  2068 => x"7451b78f",
  2069 => x"2d81f451",
  2070 => x"b48a2d80",
  2071 => x"e4b40881",
  2072 => x"2a708106",
  2073 => x"51527180",
  2074 => x"2eb33874",
  2075 => x"08852e09",
  2076 => x"8106aa38",
  2077 => x"881580f5",
  2078 => x"2d810552",
  2079 => x"71881681",
  2080 => x"b72d7181",
  2081 => x"ff068b16",
  2082 => x"80f52d54",
  2083 => x"52727227",
  2084 => x"87387288",
  2085 => x"1681b72d",
  2086 => x"7451b78f",
  2087 => x"2d80da51",
  2088 => x"b48a2d80",
  2089 => x"e4b40881",
  2090 => x"2a708106",
  2091 => x"5152718e",
  2092 => x"3880e584",
  2093 => x"08810652",
  2094 => x"80722581",
  2095 => x"c23880e5",
  2096 => x"940880e5",
  2097 => x"84088106",
  2098 => x"53538072",
  2099 => x"258438b6",
  2100 => x"a42d80e5",
  2101 => x"9c085473",
  2102 => x"802e8b38",
  2103 => x"8c13ff15",
  2104 => x"555380c1",
  2105 => x"d7047208",
  2106 => x"5271822e",
  2107 => x"a8387182",
  2108 => x"268a3871",
  2109 => x"812ead38",
  2110 => x"80c2ff04",
  2111 => x"71832eb7",
  2112 => x"3871842e",
  2113 => x"09810680",
  2114 => x"f6388813",
  2115 => x"0851b8e5",
  2116 => x"2d80c2ff",
  2117 => x"0480e59c",
  2118 => x"08518813",
  2119 => x"0852712d",
  2120 => x"80c2ff04",
  2121 => x"810b8814",
  2122 => x"082b80e2",
  2123 => x"f0083280",
  2124 => x"e2f00c80",
  2125 => x"c2d20488",
  2126 => x"1380f52d",
  2127 => x"81058b14",
  2128 => x"80f52d53",
  2129 => x"54717424",
  2130 => x"83388054",
  2131 => x"73881481",
  2132 => x"b72db7bf",
  2133 => x"2d80c2ff",
  2134 => x"04750880",
  2135 => x"2ea43875",
  2136 => x"0851b48a",
  2137 => x"2d80e4b4",
  2138 => x"08810652",
  2139 => x"71802e8c",
  2140 => x"3880e59c",
  2141 => x"08518416",
  2142 => x"0852712d",
  2143 => x"88165675",
  2144 => x"d8388054",
  2145 => x"800b80e4",
  2146 => x"c80c738f",
  2147 => x"0680e4c4",
  2148 => x"0ca05273",
  2149 => x"80e59c08",
  2150 => x"2e098106",
  2151 => x"993880e5",
  2152 => x"9808ff05",
  2153 => x"74327009",
  2154 => x"81057072",
  2155 => x"079f2a91",
  2156 => x"71315151",
  2157 => x"53537151",
  2158 => x"83842d81",
  2159 => x"14548e74",
  2160 => x"25c23880",
  2161 => x"e2f40852",
  2162 => x"7180e4b4",
  2163 => x"0c029805",
  2164 => x"0d0402f4",
  2165 => x"050dd452",
  2166 => x"81ff720c",
  2167 => x"71085381",
  2168 => x"ff720c72",
  2169 => x"882b83fe",
  2170 => x"80067208",
  2171 => x"7081ff06",
  2172 => x"51525381",
  2173 => x"ff720c72",
  2174 => x"7107882b",
  2175 => x"72087081",
  2176 => x"ff065152",
  2177 => x"5381ff72",
  2178 => x"0c727107",
  2179 => x"882b7208",
  2180 => x"7081ff06",
  2181 => x"720780e4",
  2182 => x"b40c5253",
  2183 => x"028c050d",
  2184 => x"0402f405",
  2185 => x"0d747671",
  2186 => x"81ff06d4",
  2187 => x"0c535380",
  2188 => x"e5a40885",
  2189 => x"3871892b",
  2190 => x"5271982a",
  2191 => x"d40c7190",
  2192 => x"2a7081ff",
  2193 => x"06d40c51",
  2194 => x"71882a70",
  2195 => x"81ff06d4",
  2196 => x"0c517181",
  2197 => x"ff06d40c",
  2198 => x"72902a70",
  2199 => x"81ff06d4",
  2200 => x"0c51d408",
  2201 => x"7081ff06",
  2202 => x"515182b8",
  2203 => x"bf527081",
  2204 => x"ff2e0981",
  2205 => x"06943881",
  2206 => x"ff0bd40c",
  2207 => x"d4087081",
  2208 => x"ff06ff14",
  2209 => x"54515171",
  2210 => x"e5387080",
  2211 => x"e4b40c02",
  2212 => x"8c050d04",
  2213 => x"02fc050d",
  2214 => x"81c75181",
  2215 => x"ff0bd40c",
  2216 => x"ff115170",
  2217 => x"8025f438",
  2218 => x"0284050d",
  2219 => x"0402f405",
  2220 => x"0d81ff0b",
  2221 => x"d40c9353",
  2222 => x"805287fc",
  2223 => x"80c15180",
  2224 => x"c4a12d80",
  2225 => x"e4b4088c",
  2226 => x"3881ff0b",
  2227 => x"d40c8153",
  2228 => x"80c5de04",
  2229 => x"80c5942d",
  2230 => x"ff135372",
  2231 => x"db387280",
  2232 => x"e4b40c02",
  2233 => x"8c050d04",
  2234 => x"02ec050d",
  2235 => x"810b80e5",
  2236 => x"a40c8454",
  2237 => x"d008708f",
  2238 => x"2a708106",
  2239 => x"51515372",
  2240 => x"f33872d0",
  2241 => x"0c80c594",
  2242 => x"2d80e09c",
  2243 => x"5186a02d",
  2244 => x"d008708f",
  2245 => x"2a708106",
  2246 => x"51515372",
  2247 => x"f338810b",
  2248 => x"d00cb153",
  2249 => x"805284d4",
  2250 => x"80c05180",
  2251 => x"c4a12d80",
  2252 => x"e4b40881",
  2253 => x"2e943872",
  2254 => x"822e80c4",
  2255 => x"38ff1353",
  2256 => x"72e238ff",
  2257 => x"145473ff",
  2258 => x"ab3880c5",
  2259 => x"942d83aa",
  2260 => x"52849c80",
  2261 => x"c85180c4",
  2262 => x"a12d80e4",
  2263 => x"b408812e",
  2264 => x"09810694",
  2265 => x"3880c3d2",
  2266 => x"2d80e4b4",
  2267 => x"0883ffff",
  2268 => x"06537283",
  2269 => x"aa2ea338",
  2270 => x"80c5ad2d",
  2271 => x"80c79404",
  2272 => x"80e0a851",
  2273 => x"86a02d80",
  2274 => x"5380c8f2",
  2275 => x"0480e0c0",
  2276 => x"5186a02d",
  2277 => x"805480c8",
  2278 => x"c20481ff",
  2279 => x"0bd40cb1",
  2280 => x"5480c594",
  2281 => x"2d8fcf53",
  2282 => x"805287fc",
  2283 => x"80f75180",
  2284 => x"c4a12d80",
  2285 => x"e4b40855",
  2286 => x"80e4b408",
  2287 => x"812e0981",
  2288 => x"069e3881",
  2289 => x"ff0bd40c",
  2290 => x"820a5284",
  2291 => x"9c80e951",
  2292 => x"80c4a12d",
  2293 => x"80e4b408",
  2294 => x"802e8f38",
  2295 => x"80c5942d",
  2296 => x"ff135372",
  2297 => x"c33880c8",
  2298 => x"b50481ff",
  2299 => x"0bd40c80",
  2300 => x"e4b40852",
  2301 => x"87fc80fa",
  2302 => x"5180c4a1",
  2303 => x"2d80e4b4",
  2304 => x"08b33881",
  2305 => x"ff0bd40c",
  2306 => x"d4085381",
  2307 => x"ff0bd40c",
  2308 => x"81ff0bd4",
  2309 => x"0c81ff0b",
  2310 => x"d40c81ff",
  2311 => x"0bd40c72",
  2312 => x"862a7081",
  2313 => x"06765651",
  2314 => x"53729738",
  2315 => x"80e4b408",
  2316 => x"5480c8c2",
  2317 => x"0473822e",
  2318 => x"fed338ff",
  2319 => x"145473fe",
  2320 => x"e0387380",
  2321 => x"e5a40c73",
  2322 => x"8c388152",
  2323 => x"87fc80d0",
  2324 => x"5180c4a1",
  2325 => x"2d81ff0b",
  2326 => x"d40cd008",
  2327 => x"708f2a70",
  2328 => x"81065151",
  2329 => x"5372f338",
  2330 => x"72d00c81",
  2331 => x"ff0bd40c",
  2332 => x"81537280",
  2333 => x"e4b40c02",
  2334 => x"94050d04",
  2335 => x"02e8050d",
  2336 => x"78558056",
  2337 => x"81ff0bd4",
  2338 => x"0cd00870",
  2339 => x"8f2a7081",
  2340 => x"06515153",
  2341 => x"72f33882",
  2342 => x"810bd00c",
  2343 => x"81ff0bd4",
  2344 => x"0c775287",
  2345 => x"fc80d151",
  2346 => x"80c4a12d",
  2347 => x"80dbc6df",
  2348 => x"5480e4b4",
  2349 => x"08802e8c",
  2350 => x"3880e0e0",
  2351 => x"5186a02d",
  2352 => x"80ca9a04",
  2353 => x"81ff0bd4",
  2354 => x"0cd40870",
  2355 => x"81ff0651",
  2356 => x"537281fe",
  2357 => x"2e098106",
  2358 => x"a03880ff",
  2359 => x"5380c3d2",
  2360 => x"2d80e4b4",
  2361 => x"08757084",
  2362 => x"05570cff",
  2363 => x"13537280",
  2364 => x"25eb3881",
  2365 => x"5680c9ff",
  2366 => x"04ff1454",
  2367 => x"73c63881",
  2368 => x"ff0bd40c",
  2369 => x"81ff0bd4",
  2370 => x"0cd00870",
  2371 => x"8f2a7081",
  2372 => x"06515153",
  2373 => x"72f33872",
  2374 => x"d00c7580",
  2375 => x"e4b40c02",
  2376 => x"98050d04",
  2377 => x"02e8050d",
  2378 => x"77797b58",
  2379 => x"55558053",
  2380 => x"727625a5",
  2381 => x"38747081",
  2382 => x"055680f5",
  2383 => x"2d747081",
  2384 => x"055680f5",
  2385 => x"2d525271",
  2386 => x"712e8738",
  2387 => x"815180ca",
  2388 => x"db048113",
  2389 => x"5380cab0",
  2390 => x"04805170",
  2391 => x"80e4b40c",
  2392 => x"0298050d",
  2393 => x"0402ec05",
  2394 => x"0d765574",
  2395 => x"802e80c4",
  2396 => x"389a1580",
  2397 => x"e02d5180",
  2398 => x"d9a02d80",
  2399 => x"e4b40880",
  2400 => x"e4b40880",
  2401 => x"ebd80c80",
  2402 => x"e4b40854",
  2403 => x"5480ebb4",
  2404 => x"08802e9b",
  2405 => x"38941580",
  2406 => x"e02d5180",
  2407 => x"d9a02d80",
  2408 => x"e4b40890",
  2409 => x"2b83fff0",
  2410 => x"0a067075",
  2411 => x"07515372",
  2412 => x"80ebd80c",
  2413 => x"80ebd808",
  2414 => x"5372802e",
  2415 => x"9e3880eb",
  2416 => x"ac08fe14",
  2417 => x"712980eb",
  2418 => x"c0080580",
  2419 => x"ebdc0c70",
  2420 => x"842b80eb",
  2421 => x"b80c5480",
  2422 => x"cc8a0480",
  2423 => x"ebc40880",
  2424 => x"ebd80c80",
  2425 => x"ebc80880",
  2426 => x"ebdc0c80",
  2427 => x"ebb40880",
  2428 => x"2e8c3880",
  2429 => x"ebac0884",
  2430 => x"2b5380cc",
  2431 => x"850480eb",
  2432 => x"cc08842b",
  2433 => x"537280eb",
  2434 => x"b80c0294",
  2435 => x"050d0402",
  2436 => x"d8050d80",
  2437 => x"0b80ebb4",
  2438 => x"0c845480",
  2439 => x"c5e82d80",
  2440 => x"e4b40880",
  2441 => x"2e993880",
  2442 => x"e5a85280",
  2443 => x"5180c8fc",
  2444 => x"2d80e4b4",
  2445 => x"08802e87",
  2446 => x"38fe5480",
  2447 => x"ccc704ff",
  2448 => x"14547380",
  2449 => x"24d53873",
  2450 => x"8e3880e0",
  2451 => x"f05186a0",
  2452 => x"2d735580",
  2453 => x"d2ab0480",
  2454 => x"56810b80",
  2455 => x"ebe00c88",
  2456 => x"5380e184",
  2457 => x"5280e5de",
  2458 => x"5180caa4",
  2459 => x"2d80e4b4",
  2460 => x"08762e09",
  2461 => x"81068938",
  2462 => x"80e4b408",
  2463 => x"80ebe00c",
  2464 => x"885380e1",
  2465 => x"905280e5",
  2466 => x"fa5180ca",
  2467 => x"a42d80e4",
  2468 => x"b4088938",
  2469 => x"80e4b408",
  2470 => x"80ebe00c",
  2471 => x"80ebe008",
  2472 => x"802e8185",
  2473 => x"3880e8ee",
  2474 => x"0b80f52d",
  2475 => x"80e8ef0b",
  2476 => x"80f52d71",
  2477 => x"982b7190",
  2478 => x"2b0780e8",
  2479 => x"f00b80f5",
  2480 => x"2d70882b",
  2481 => x"720780e8",
  2482 => x"f10b80f5",
  2483 => x"2d710780",
  2484 => x"e9a60b80",
  2485 => x"f52d80e9",
  2486 => x"a70b80f5",
  2487 => x"2d71882b",
  2488 => x"07535f54",
  2489 => x"525a5657",
  2490 => x"557381ab",
  2491 => x"aa2e0981",
  2492 => x"06903875",
  2493 => x"5180d8ef",
  2494 => x"2d80e4b4",
  2495 => x"085680ce",
  2496 => x"91047382",
  2497 => x"d4d52e89",
  2498 => x"3880e19c",
  2499 => x"5180cee1",
  2500 => x"0480e5a8",
  2501 => x"52755180",
  2502 => x"c8fc2d80",
  2503 => x"e4b40855",
  2504 => x"80e4b408",
  2505 => x"802e8483",
  2506 => x"38885380",
  2507 => x"e1905280",
  2508 => x"e5fa5180",
  2509 => x"caa42d80",
  2510 => x"e4b4088b",
  2511 => x"38810b80",
  2512 => x"ebb40c80",
  2513 => x"cee80488",
  2514 => x"5380e184",
  2515 => x"5280e5de",
  2516 => x"5180caa4",
  2517 => x"2d80e4b4",
  2518 => x"08802e8c",
  2519 => x"3880e1b0",
  2520 => x"5186a02d",
  2521 => x"80cfc704",
  2522 => x"80e9a60b",
  2523 => x"80f52d54",
  2524 => x"7380d52e",
  2525 => x"09810680",
  2526 => x"ce3880e9",
  2527 => x"a70b80f5",
  2528 => x"2d547381",
  2529 => x"aa2e0981",
  2530 => x"06bd3880",
  2531 => x"0b80e5a8",
  2532 => x"0b80f52d",
  2533 => x"56547481",
  2534 => x"e92e8338",
  2535 => x"81547481",
  2536 => x"eb2e8c38",
  2537 => x"80557375",
  2538 => x"2e098106",
  2539 => x"82fd3880",
  2540 => x"e5b30b80",
  2541 => x"f52d5574",
  2542 => x"8e3880e5",
  2543 => x"b40b80f5",
  2544 => x"2d547382",
  2545 => x"2e873880",
  2546 => x"5580d2ab",
  2547 => x"0480e5b5",
  2548 => x"0b80f52d",
  2549 => x"7080ebac",
  2550 => x"0cff0580",
  2551 => x"ebb00c80",
  2552 => x"e5b60b80",
  2553 => x"f52d80e5",
  2554 => x"b70b80f5",
  2555 => x"2d587605",
  2556 => x"77828029",
  2557 => x"057080eb",
  2558 => x"bc0c80e5",
  2559 => x"b80b80f5",
  2560 => x"2d7080eb",
  2561 => x"d00c80eb",
  2562 => x"b4085957",
  2563 => x"5876802e",
  2564 => x"81b93888",
  2565 => x"5380e190",
  2566 => x"5280e5fa",
  2567 => x"5180caa4",
  2568 => x"2d80e4b4",
  2569 => x"08828438",
  2570 => x"80ebac08",
  2571 => x"70842b80",
  2572 => x"ebb80c70",
  2573 => x"80ebcc0c",
  2574 => x"80e5cd0b",
  2575 => x"80f52d80",
  2576 => x"e5cc0b80",
  2577 => x"f52d7182",
  2578 => x"80290580",
  2579 => x"e5ce0b80",
  2580 => x"f52d7084",
  2581 => x"80802912",
  2582 => x"80e5cf0b",
  2583 => x"80f52d70",
  2584 => x"81800a29",
  2585 => x"127080eb",
  2586 => x"d40c80eb",
  2587 => x"d0087129",
  2588 => x"80ebbc08",
  2589 => x"057080eb",
  2590 => x"c00c80e5",
  2591 => x"d50b80f5",
  2592 => x"2d80e5d4",
  2593 => x"0b80f52d",
  2594 => x"71828029",
  2595 => x"0580e5d6",
  2596 => x"0b80f52d",
  2597 => x"70848080",
  2598 => x"291280e5",
  2599 => x"d70b80f5",
  2600 => x"2d70982b",
  2601 => x"81f00a06",
  2602 => x"72057080",
  2603 => x"ebc40cfe",
  2604 => x"117e2977",
  2605 => x"0580ebc8",
  2606 => x"0c525952",
  2607 => x"43545e51",
  2608 => x"5259525d",
  2609 => x"57595780",
  2610 => x"d2a30480",
  2611 => x"e5ba0b80",
  2612 => x"f52d80e5",
  2613 => x"b90b80f5",
  2614 => x"2d718280",
  2615 => x"29057080",
  2616 => x"ebb80c70",
  2617 => x"a02983ff",
  2618 => x"0570892a",
  2619 => x"7080ebcc",
  2620 => x"0c80e5bf",
  2621 => x"0b80f52d",
  2622 => x"80e5be0b",
  2623 => x"80f52d71",
  2624 => x"82802905",
  2625 => x"7080ebd4",
  2626 => x"0c7b7129",
  2627 => x"1e7080eb",
  2628 => x"c80c7d80",
  2629 => x"ebc40c73",
  2630 => x"0580ebc0",
  2631 => x"0c555e51",
  2632 => x"51555580",
  2633 => x"5180cae5",
  2634 => x"2d815574",
  2635 => x"80e4b40c",
  2636 => x"02a8050d",
  2637 => x"0402ec05",
  2638 => x"0d767087",
  2639 => x"2c7180ff",
  2640 => x"06555654",
  2641 => x"80ebb408",
  2642 => x"8a387388",
  2643 => x"2c7481ff",
  2644 => x"06545580",
  2645 => x"e5a85280",
  2646 => x"ebbc0815",
  2647 => x"5180c8fc",
  2648 => x"2d80e4b4",
  2649 => x"085480e4",
  2650 => x"b408802e",
  2651 => x"bb3880eb",
  2652 => x"b408802e",
  2653 => x"9c387284",
  2654 => x"2980e5a8",
  2655 => x"05700852",
  2656 => x"5380d8ef",
  2657 => x"2d80e4b4",
  2658 => x"08f00a06",
  2659 => x"5380d3a6",
  2660 => x"04721080",
  2661 => x"e5a80570",
  2662 => x"80e02d52",
  2663 => x"5380d9a0",
  2664 => x"2d80e4b4",
  2665 => x"08537254",
  2666 => x"7380e4b4",
  2667 => x"0c029405",
  2668 => x"0d0402e0",
  2669 => x"050d7970",
  2670 => x"842c80eb",
  2671 => x"dc080571",
  2672 => x"8f065255",
  2673 => x"53728b38",
  2674 => x"80e5a852",
  2675 => x"735180c8",
  2676 => x"fc2d72a0",
  2677 => x"2980e5a8",
  2678 => x"05548074",
  2679 => x"80f52d56",
  2680 => x"5374732e",
  2681 => x"83388153",
  2682 => x"7481e52e",
  2683 => x"81f53881",
  2684 => x"70740654",
  2685 => x"5872802e",
  2686 => x"81e9388b",
  2687 => x"1480f52d",
  2688 => x"70832a79",
  2689 => x"06585676",
  2690 => x"9c3880e2",
  2691 => x"f8085372",
  2692 => x"89387280",
  2693 => x"e9a80b81",
  2694 => x"b72d7680",
  2695 => x"e2f80c73",
  2696 => x"5380d5e5",
  2697 => x"04758f2e",
  2698 => x"09810681",
  2699 => x"b638749f",
  2700 => x"068d2980",
  2701 => x"e99b1151",
  2702 => x"53811480",
  2703 => x"f52d7370",
  2704 => x"81055581",
  2705 => x"b72d8314",
  2706 => x"80f52d73",
  2707 => x"70810555",
  2708 => x"81b72d85",
  2709 => x"1480f52d",
  2710 => x"73708105",
  2711 => x"5581b72d",
  2712 => x"871480f5",
  2713 => x"2d737081",
  2714 => x"055581b7",
  2715 => x"2d891480",
  2716 => x"f52d7370",
  2717 => x"81055581",
  2718 => x"b72d8e14",
  2719 => x"80f52d73",
  2720 => x"70810555",
  2721 => x"81b72d90",
  2722 => x"1480f52d",
  2723 => x"73708105",
  2724 => x"5581b72d",
  2725 => x"921480f5",
  2726 => x"2d737081",
  2727 => x"055581b7",
  2728 => x"2d941480",
  2729 => x"f52d7370",
  2730 => x"81055581",
  2731 => x"b72d9614",
  2732 => x"80f52d73",
  2733 => x"70810555",
  2734 => x"81b72d98",
  2735 => x"1480f52d",
  2736 => x"73708105",
  2737 => x"5581b72d",
  2738 => x"9c1480f5",
  2739 => x"2d737081",
  2740 => x"055581b7",
  2741 => x"2d9e1480",
  2742 => x"f52d7381",
  2743 => x"b72d7780",
  2744 => x"e2f80c80",
  2745 => x"537280e4",
  2746 => x"b40c02a0",
  2747 => x"050d0402",
  2748 => x"cc050d7e",
  2749 => x"605e5a80",
  2750 => x"0b80ebd8",
  2751 => x"0880ebdc",
  2752 => x"08595c56",
  2753 => x"805880eb",
  2754 => x"b808782e",
  2755 => x"81be3877",
  2756 => x"8f06a017",
  2757 => x"57547392",
  2758 => x"3880e5a8",
  2759 => x"52765181",
  2760 => x"175780c8",
  2761 => x"fc2d80e5",
  2762 => x"a8568076",
  2763 => x"80f52d56",
  2764 => x"5474742e",
  2765 => x"83388154",
  2766 => x"7481e52e",
  2767 => x"81823881",
  2768 => x"70750655",
  2769 => x"5c73802e",
  2770 => x"80f6388b",
  2771 => x"1680f52d",
  2772 => x"98065978",
  2773 => x"80ea388b",
  2774 => x"537c5275",
  2775 => x"5180caa4",
  2776 => x"2d80e4b4",
  2777 => x"0880d938",
  2778 => x"9c160851",
  2779 => x"80d8ef2d",
  2780 => x"80e4b408",
  2781 => x"841b0c9a",
  2782 => x"1680e02d",
  2783 => x"5180d9a0",
  2784 => x"2d80e4b4",
  2785 => x"0880e4b4",
  2786 => x"08881c0c",
  2787 => x"80e4b408",
  2788 => x"555580eb",
  2789 => x"b408802e",
  2790 => x"9a389416",
  2791 => x"80e02d51",
  2792 => x"80d9a02d",
  2793 => x"80e4b408",
  2794 => x"902b83ff",
  2795 => x"f00a0670",
  2796 => x"16515473",
  2797 => x"881b0c78",
  2798 => x"7a0c7b54",
  2799 => x"80d88a04",
  2800 => x"81185880",
  2801 => x"ebb80878",
  2802 => x"26fec438",
  2803 => x"80ebb408",
  2804 => x"802eb538",
  2805 => x"7a5180d2",
  2806 => x"b52d80e4",
  2807 => x"b40880e4",
  2808 => x"b40880ff",
  2809 => x"fffff806",
  2810 => x"555b7380",
  2811 => x"fffffff8",
  2812 => x"2e963880",
  2813 => x"e4b408fe",
  2814 => x"0580ebac",
  2815 => x"082980eb",
  2816 => x"c0080557",
  2817 => x"80d68404",
  2818 => x"80547380",
  2819 => x"e4b40c02",
  2820 => x"b4050d04",
  2821 => x"02f4050d",
  2822 => x"74700881",
  2823 => x"05710c70",
  2824 => x"0880ebb0",
  2825 => x"08065353",
  2826 => x"71903888",
  2827 => x"13085180",
  2828 => x"d2b52d80",
  2829 => x"e4b40888",
  2830 => x"140c810b",
  2831 => x"80e4b40c",
  2832 => x"028c050d",
  2833 => x"0402f005",
  2834 => x"0d758811",
  2835 => x"08fe0580",
  2836 => x"ebac0829",
  2837 => x"80ebc008",
  2838 => x"11720880",
  2839 => x"ebb00806",
  2840 => x"05795553",
  2841 => x"545480c8",
  2842 => x"fc2d0290",
  2843 => x"050d0402",
  2844 => x"f4050d74",
  2845 => x"70882a83",
  2846 => x"fe800670",
  2847 => x"72982a07",
  2848 => x"72882b87",
  2849 => x"fc808006",
  2850 => x"73982b81",
  2851 => x"f00a0671",
  2852 => x"73070780",
  2853 => x"e4b40c56",
  2854 => x"51535102",
  2855 => x"8c050d04",
  2856 => x"02f8050d",
  2857 => x"028e0580",
  2858 => x"f52d7488",
  2859 => x"2b077083",
  2860 => x"ffff0680",
  2861 => x"e4b40c51",
  2862 => x"0288050d",
  2863 => x"0402f405",
  2864 => x"0d747678",
  2865 => x"53545280",
  2866 => x"71259738",
  2867 => x"72708105",
  2868 => x"5480f52d",
  2869 => x"72708105",
  2870 => x"5481b72d",
  2871 => x"ff115170",
  2872 => x"eb388072",
  2873 => x"81b72d02",
  2874 => x"8c050d04",
  2875 => x"02e8050d",
  2876 => x"77568070",
  2877 => x"56547376",
  2878 => x"24b73880",
  2879 => x"ebb80874",
  2880 => x"2eaf3873",
  2881 => x"5180d3b2",
  2882 => x"2d80e4b4",
  2883 => x"0880e4b4",
  2884 => x"08098105",
  2885 => x"7080e4b4",
  2886 => x"08079f2a",
  2887 => x"77058117",
  2888 => x"57575353",
  2889 => x"74762489",
  2890 => x"3880ebb8",
  2891 => x"087426d3",
  2892 => x"387280e4",
  2893 => x"b40c0298",
  2894 => x"050d0402",
  2895 => x"f0050d80",
  2896 => x"e4b00816",
  2897 => x"5180d9ec",
  2898 => x"2d80e4b4",
  2899 => x"08802ea0",
  2900 => x"388b5380",
  2901 => x"e4b40852",
  2902 => x"80e9a851",
  2903 => x"80d9bd2d",
  2904 => x"80ebe408",
  2905 => x"5473802e",
  2906 => x"873880e9",
  2907 => x"a851732d",
  2908 => x"0290050d",
  2909 => x"0402dc05",
  2910 => x"0d80705a",
  2911 => x"557480e4",
  2912 => x"b00825b5",
  2913 => x"3880ebb8",
  2914 => x"08752ead",
  2915 => x"38785180",
  2916 => x"d3b22d80",
  2917 => x"e4b40809",
  2918 => x"81057080",
  2919 => x"e4b40807",
  2920 => x"9f2a7605",
  2921 => x"811b5b56",
  2922 => x"547480e4",
  2923 => x"b0082589",
  2924 => x"3880ebb8",
  2925 => x"087926d5",
  2926 => x"38805578",
  2927 => x"80ebb808",
  2928 => x"2781e438",
  2929 => x"785180d3",
  2930 => x"b22d80e4",
  2931 => x"b408802e",
  2932 => x"81b43880",
  2933 => x"e4b4088b",
  2934 => x"0580f52d",
  2935 => x"70842a70",
  2936 => x"81067710",
  2937 => x"78842b80",
  2938 => x"e9a80b80",
  2939 => x"f52d5c5c",
  2940 => x"53515556",
  2941 => x"73802e80",
  2942 => x"ce387416",
  2943 => x"822b80dd",
  2944 => x"cb0b80e3",
  2945 => x"84120c54",
  2946 => x"77753110",
  2947 => x"80ebe811",
  2948 => x"55569074",
  2949 => x"70810556",
  2950 => x"81b72da0",
  2951 => x"7481b72d",
  2952 => x"7681ff06",
  2953 => x"81165854",
  2954 => x"73802e8b",
  2955 => x"389c5380",
  2956 => x"e9a85280",
  2957 => x"dcbe048b",
  2958 => x"5380e4b4",
  2959 => x"085280eb",
  2960 => x"ea165180",
  2961 => x"dcfc0474",
  2962 => x"16822b80",
  2963 => x"dabb0b80",
  2964 => x"e384120c",
  2965 => x"547681ff",
  2966 => x"06811658",
  2967 => x"5473802e",
  2968 => x"8b389c53",
  2969 => x"80e9a852",
  2970 => x"80dcf304",
  2971 => x"8b5380e4",
  2972 => x"b4085277",
  2973 => x"75311080",
  2974 => x"ebe80551",
  2975 => x"765580d9",
  2976 => x"bd2d80dd",
  2977 => x"9b047490",
  2978 => x"29753170",
  2979 => x"1080ebe8",
  2980 => x"05515480",
  2981 => x"e4b40874",
  2982 => x"81b72d81",
  2983 => x"1959748b",
  2984 => x"24a43880",
  2985 => x"dbbb0474",
  2986 => x"90297531",
  2987 => x"701080eb",
  2988 => x"e8058c77",
  2989 => x"31575154",
  2990 => x"807481b7",
  2991 => x"2d9e14ff",
  2992 => x"16565474",
  2993 => x"f33802a4",
  2994 => x"050d0402",
  2995 => x"fc050d80",
  2996 => x"e4b00813",
  2997 => x"5180d9ec",
  2998 => x"2d80e4b4",
  2999 => x"08802e8a",
  3000 => x"3880e4b4",
  3001 => x"085180ca",
  3002 => x"e52d800b",
  3003 => x"80e4b00c",
  3004 => x"80daf52d",
  3005 => x"b7bf2d02",
  3006 => x"84050d04",
  3007 => x"02fc050d",
  3008 => x"725170fd",
  3009 => x"2eb23870",
  3010 => x"fd248b38",
  3011 => x"70fc2e80",
  3012 => x"d03880de",
  3013 => x"eb0470fe",
  3014 => x"2eb93870",
  3015 => x"ff2e0981",
  3016 => x"0680c838",
  3017 => x"80e4b008",
  3018 => x"5170802e",
  3019 => x"be38ff11",
  3020 => x"80e4b00c",
  3021 => x"80deeb04",
  3022 => x"80e4b008",
  3023 => x"f0057080",
  3024 => x"e4b00c51",
  3025 => x"708025a3",
  3026 => x"38800b80",
  3027 => x"e4b00c80",
  3028 => x"deeb0480",
  3029 => x"e4b00881",
  3030 => x"0580e4b0",
  3031 => x"0c80deeb",
  3032 => x"0480e4b0",
  3033 => x"08900580",
  3034 => x"e4b00c80",
  3035 => x"daf52db7",
  3036 => x"bf2d0284",
  3037 => x"050d0402",
  3038 => x"fc050d80",
  3039 => x"0b80e4b0",
  3040 => x"0c80daf5",
  3041 => x"2db6bb2d",
  3042 => x"80e4b408",
  3043 => x"80e4a00c",
  3044 => x"80e2fc51",
  3045 => x"b8e52d02",
  3046 => x"84050d04",
  3047 => x"7180ebe4",
  3048 => x"0c040000",
  3049 => x"00ffffff",
  3050 => x"ff00ffff",
  3051 => x"ffff00ff",
  3052 => x"ffffff00",
  3053 => x"52657365",
  3054 => x"74204e45",
  3055 => x"53000000",
  3056 => x"5363616e",
  3057 => x"6c696e65",
  3058 => x"73000000",
  3059 => x"4c6f6164",
  3060 => x"20524f4d",
  3061 => x"20100000",
  3062 => x"45786974",
  3063 => x"00000000",
  3064 => x"524f4d20",
  3065 => x"6c6f6164",
  3066 => x"696e6720",
  3067 => x"6661696c",
  3068 => x"65640000",
  3069 => x"4f4b0000",
  3070 => x"496e6974",
  3071 => x"69616c69",
  3072 => x"7a696e67",
  3073 => x"20534420",
  3074 => x"63617264",
  3075 => x"0a000000",
  3076 => x"16200000",
  3077 => x"14200000",
  3078 => x"15200000",
  3079 => x"53442069",
  3080 => x"6e69742e",
  3081 => x"2e2e0a00",
  3082 => x"53442063",
  3083 => x"61726420",
  3084 => x"72657365",
  3085 => x"74206661",
  3086 => x"696c6564",
  3087 => x"210a0000",
  3088 => x"53444843",
  3089 => x"20657272",
  3090 => x"6f72210a",
  3091 => x"00000000",
  3092 => x"57726974",
  3093 => x"65206661",
  3094 => x"696c6564",
  3095 => x"0a000000",
  3096 => x"52656164",
  3097 => x"20666169",
  3098 => x"6c65640a",
  3099 => x"00000000",
  3100 => x"43617264",
  3101 => x"20696e69",
  3102 => x"74206661",
  3103 => x"696c6564",
  3104 => x"0a000000",
  3105 => x"46415431",
  3106 => x"36202020",
  3107 => x"00000000",
  3108 => x"46415433",
  3109 => x"32202020",
  3110 => x"00000000",
  3111 => x"4e6f2070",
  3112 => x"61727469",
  3113 => x"74696f6e",
  3114 => x"20736967",
  3115 => x"0a000000",
  3116 => x"42616420",
  3117 => x"70617274",
  3118 => x"0a000000",
  3119 => x"4261636b",
  3120 => x"00000000",
  3121 => x"00000002",
  3122 => x"00000002",
  3123 => x"00002fb4",
  3124 => x"0000035a",
  3125 => x"00000001",
  3126 => x"00002fc0",
  3127 => x"00000000",
  3128 => x"00000002",
  3129 => x"00002fcc",
  3130 => x"00002f77",
  3131 => x"00000002",
  3132 => x"00002fd8",
  3133 => x"00001b58",
  3134 => x"00000000",
  3135 => x"00000000",
  3136 => x"00000000",
  3137 => x"00000004",
  3138 => x"00002fe0",
  3139 => x"00003104",
  3140 => x"00000004",
  3141 => x"00002ff4",
  3142 => x"000030c8",
  3143 => x"00000000",
  3144 => x"00000000",
  3145 => x"00000000",
  3146 => x"00000000",
  3147 => x"00000000",
  3148 => x"00000000",
  3149 => x"00000000",
  3150 => x"00000000",
  3151 => x"00000000",
  3152 => x"00000000",
  3153 => x"00000000",
  3154 => x"00000000",
  3155 => x"00000000",
  3156 => x"00000000",
  3157 => x"00000000",
  3158 => x"00000000",
  3159 => x"00000000",
  3160 => x"00000000",
  3161 => x"00000000",
  3162 => x"00000000",
  3163 => x"00000000",
  3164 => x"00000000",
  3165 => x"00000000",
  3166 => x"00000000",
  3167 => x"00000002",
  3168 => x"000035e8",
  3169 => x"00002d3b",
  3170 => x"00000002",
  3171 => x"00003606",
  3172 => x"00002d3b",
  3173 => x"00000002",
  3174 => x"00003624",
  3175 => x"00002d3b",
  3176 => x"00000002",
  3177 => x"00003642",
  3178 => x"00002d3b",
  3179 => x"00000002",
  3180 => x"00003660",
  3181 => x"00002d3b",
  3182 => x"00000002",
  3183 => x"0000367e",
  3184 => x"00002d3b",
  3185 => x"00000002",
  3186 => x"0000369c",
  3187 => x"00002d3b",
  3188 => x"00000002",
  3189 => x"000036ba",
  3190 => x"00002d3b",
  3191 => x"00000002",
  3192 => x"000036d8",
  3193 => x"00002d3b",
  3194 => x"00000002",
  3195 => x"000036f6",
  3196 => x"00002d3b",
  3197 => x"00000002",
  3198 => x"00003714",
  3199 => x"00002d3b",
  3200 => x"00000002",
  3201 => x"00003732",
  3202 => x"00002d3b",
  3203 => x"00000002",
  3204 => x"00003750",
  3205 => x"00002d3b",
  3206 => x"00000004",
  3207 => x"000030bc",
  3208 => x"00000000",
  3209 => x"00000000",
  3210 => x"00000000",
  3211 => x"00002efc",
  3212 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

