-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;


entity bootrom is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of bootrom is


  type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"F3",x"ED",x"56",x"C3",x"80",x"00",x"FF",x"FF", -- 0x0000
    x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0008
    x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0010
    x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0018
    x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0020
    x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0028
    x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0030
    x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0038
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0040
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0048
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0050
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"ED",x"45", -- 0x0060
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0068
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0070
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0078
    x"31",x"FF",x"FF",x"CD",x"00",x"22",x"CD",x"99", -- 0x0080
    x"02",x"C3",x"00",x"01",x"FF",x"FF",x"FF",x"FF", -- 0x0088
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0090
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0098
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00F8
    x"76",x"18",x"FD",x"CD",x"05",x"1E",x"21",x"01", -- 0x0100
    x"0A",x"E5",x"CD",x"2A",x"1E",x"21",x"45",x"01", -- 0x0108
    x"E3",x"CD",x"B4",x"1F",x"F1",x"C1",x"E1",x"E5", -- 0x0110
    x"C5",x"E5",x"CD",x"B4",x"1F",x"21",x"01",x"0C", -- 0x0118
    x"E3",x"CD",x"2A",x"1E",x"21",x"4D",x"01",x"E3", -- 0x0120
    x"CD",x"B4",x"1F",x"F1",x"3E",x"FF",x"D3",x"E7", -- 0x0128
    x"3E",x"02",x"D3",x"FE",x"18",x"FE",x"5C",x"7C", -- 0x0130
    x"2F",x"2D",x"00",x"06",x"04",x"05",x"03",x"AB", -- 0x0138
    x"0B",x"01",x"02",x"C7",x"D8",x"45",x"72",x"72", -- 0x0140
    x"6F",x"72",x"3A",x"20",x"00",x"50",x"72",x"65", -- 0x0148
    x"73",x"73",x"20",x"62",x"75",x"74",x"74",x"6F", -- 0x0150
    x"6E",x"20",x"31",x"20",x"74",x"6F",x"20",x"74", -- 0x0158
    x"72",x"79",x"20",x"61",x"67",x"61",x"69",x"6E", -- 0x0160
    x"00",x"01",x"00",x"00",x"21",x"02",x"00",x"39", -- 0x0168
    x"79",x"96",x"78",x"23",x"9E",x"E2",x"7A",x"01", -- 0x0170
    x"EE",x"80",x"F0",x"00",x"03",x"18",x"ED",x"FD", -- 0x0178
    x"21",x"02",x"00",x"FD",x"39",x"FD",x"7E",x"00", -- 0x0180
    x"E6",x"F0",x"07",x"07",x"07",x"07",x"E6",x"0F", -- 0x0188
    x"4F",x"FD",x"7E",x"00",x"E6",x"0F",x"07",x"07", -- 0x0190
    x"07",x"07",x"E6",x"F0",x"B1",x"FD",x"77",x"00", -- 0x0198
    x"FD",x"7E",x"00",x"E6",x"CC",x"4F",x"CB",x"39", -- 0x01A0
    x"CB",x"39",x"FD",x"7E",x"00",x"E6",x"33",x"87", -- 0x01A8
    x"87",x"B1",x"FD",x"77",x"00",x"FD",x"7E",x"00", -- 0x01B0
    x"E6",x"AA",x"4F",x"CB",x"39",x"FD",x"7E",x"00", -- 0x01B8
    x"E6",x"55",x"87",x"B1",x"FD",x"77",x"00",x"FD", -- 0x01C0
    x"6E",x"00",x"C9",x"21",x"42",x"01",x"4E",x"21", -- 0x01C8
    x"02",x"F8",x"71",x"F5",x"FD",x"21",x"28",x"FA", -- 0x01D0
    x"FD",x"5E",x"00",x"FD",x"56",x"01",x"FD",x"4E", -- 0x01D8
    x"02",x"FD",x"6E",x"03",x"F1",x"06",x"10",x"CB", -- 0x01E0
    x"3D",x"CB",x"19",x"CB",x"1A",x"CB",x"1B",x"10", -- 0x01E8
    x"F6",x"21",x"03",x"F8",x"73",x"F5",x"FD",x"5E", -- 0x01F0
    x"00",x"FD",x"56",x"01",x"FD",x"4E",x"02",x"FD", -- 0x01F8
    x"6E",x"03",x"F1",x"06",x"08",x"CB",x"3D",x"CB", -- 0x0200
    x"19",x"CB",x"1A",x"CB",x"1B",x"10",x"F6",x"21", -- 0x0208
    x"04",x"F8",x"73",x"FD",x"4E",x"00",x"21",x"05", -- 0x0210
    x"F8",x"71",x"01",x"00",x"00",x"59",x"50",x"FD", -- 0x0218
    x"21",x"02",x"00",x"FD",x"39",x"FD",x"7E",x"00", -- 0x0220
    x"83",x"5F",x"FD",x"7E",x"01",x"8A",x"57",x"1A", -- 0x0228
    x"57",x"21",x"04",x"00",x"09",x"3E",x"02",x"85", -- 0x0230
    x"6F",x"3E",x"F8",x"8C",x"67",x"E5",x"C5",x"D5", -- 0x0238
    x"33",x"CD",x"7F",x"01",x"33",x"5D",x"C1",x"E1", -- 0x0240
    x"73",x"03",x"78",x"EE",x"80",x"D6",x"81",x"38", -- 0x0248
    x"CC",x"21",x"3B",x"01",x"46",x"C5",x"33",x"CD", -- 0x0250
    x"F5",x"08",x"33",x"21",x"02",x"F8",x"E5",x"CD", -- 0x0258
    x"23",x"09",x"F1",x"01",x"36",x"01",x"2A",x"65", -- 0x0260
    x"FC",x"26",x"00",x"09",x"46",x"C5",x"33",x"CD", -- 0x0268
    x"4B",x"1E",x"33",x"3E",x"08",x"F5",x"33",x"CD", -- 0x0270
    x"4B",x"1E",x"33",x"FD",x"21",x"65",x"FC",x"FD", -- 0x0278
    x"7E",x"00",x"3C",x"E6",x"03",x"FD",x"77",x"00", -- 0x0280
    x"21",x"3D",x"01",x"46",x"C5",x"33",x"CD",x"0A", -- 0x0288
    x"09",x"33",x"7D",x"E6",x"01",x"3D",x"28",x"F0", -- 0x0290
    x"C9",x"21",x"E8",x"FF",x"39",x"F9",x"21",x"00", -- 0x0298
    x"60",x"E3",x"21",x"02",x"F8",x"36",x"00",x"5D", -- 0x02A0
    x"54",x"13",x"01",x"25",x"02",x"ED",x"B0",x"3E", -- 0x02A8
    x"00",x"01",x"3B",x"24",x"ED",x"79",x"3E",x"25", -- 0x02B0
    x"DB",x"3B",x"3E",x"01",x"01",x"3B",x"24",x"ED", -- 0x02B8
    x"79",x"3E",x"25",x"DB",x"3B",x"3E",x"02",x"01", -- 0x02C0
    x"3B",x"24",x"ED",x"79",x"3E",x"25",x"DB",x"3B", -- 0x02C8
    x"3E",x"10",x"01",x"3B",x"24",x"ED",x"79",x"3E", -- 0x02D0
    x"25",x"DB",x"3B",x"CD",x"05",x"1E",x"3E",x"01", -- 0x02D8
    x"D3",x"FE",x"21",x"04",x"04",x"E5",x"CD",x"2A", -- 0x02E0
    x"1E",x"21",x"2A",x"06",x"E3",x"CD",x"B4",x"1F", -- 0x02E8
    x"21",x"0B",x"08",x"E3",x"CD",x"2A",x"1E",x"21", -- 0x02F0
    x"43",x"06",x"E3",x"CD",x"B4",x"1F",x"21",x"02", -- 0x02F8
    x"0A",x"E3",x"CD",x"2A",x"1E",x"21",x"4E",x"06", -- 0x0300
    x"E3",x"CD",x"B4",x"1F",x"21",x"05",x"0C",x"E3", -- 0x0308
    x"CD",x"2A",x"1E",x"21",x"6B",x"06",x"E3",x"CD", -- 0x0310
    x"B4",x"1F",x"21",x"19",x"17",x"E3",x"CD",x"2A", -- 0x0318
    x"1E",x"21",x"82",x"06",x"E3",x"CD",x"B4",x"1F", -- 0x0320
    x"F1",x"3E",x"BF",x"DB",x"FE",x"E6",x"01",x"3D", -- 0x0328
    x"28",x"F7",x"21",x"07",x"0F",x"E5",x"CD",x"2A", -- 0x0330
    x"1E",x"21",x"89",x"06",x"E3",x"CD",x"B4",x"1F", -- 0x0338
    x"F1",x"3E",x"DF",x"DB",x"FE",x"E6",x"10",x"07", -- 0x0340
    x"07",x"07",x"07",x"E6",x"0F",x"3D",x"28",x"F1", -- 0x0348
    x"CD",x"05",x"1E",x"3E",x"01",x"01",x"3B",x"30", -- 0x0350
    x"ED",x"79",x"21",x"00",x"F8",x"36",x"0A",x"3A", -- 0x0358
    x"00",x"F8",x"B7",x"28",x"28",x"CD",x"6A",x"07", -- 0x0360
    x"7D",x"B7",x"20",x"08",x"21",x"9D",x"06",x"E5", -- 0x0368
    x"CD",x"03",x"01",x"F1",x"CD",x"5E",x"0D",x"7D", -- 0x0370
    x"B7",x"20",x"12",x"21",x"00",x"F8",x"35",x"01", -- 0x0378
    x"E8",x"FD",x"59",x"50",x"1B",x"4B",x"7A",x"47", -- 0x0380
    x"B3",x"20",x"F7",x"18",x"D2",x"3A",x"00",x"F8", -- 0x0388
    x"B7",x"20",x"08",x"21",x"B6",x"06",x"E5",x"CD", -- 0x0390
    x"03",x"01",x"F1",x"21",x"06",x"00",x"39",x"FD", -- 0x0398
    x"21",x"12",x"00",x"FD",x"39",x"FD",x"75",x"00", -- 0x03A0
    x"FD",x"74",x"01",x"FD",x"4E",x"00",x"FD",x"46", -- 0x03A8
    x"01",x"2A",x"63",x"FC",x"E5",x"C5",x"CD",x"BE", -- 0x03B0
    x"15",x"F1",x"F1",x"7D",x"B7",x"20",x"08",x"21", -- 0x03B8
    x"D0",x"06",x"E5",x"CD",x"03",x"01",x"F1",x"21", -- 0x03C0
    x"12",x"00",x"39",x"7E",x"23",x"66",x"6F",x"11", -- 0x03C8
    x"04",x"00",x"19",x"7E",x"FD",x"21",x"14",x"00", -- 0x03D0
    x"FD",x"39",x"FD",x"77",x"00",x"23",x"7E",x"FD", -- 0x03D8
    x"77",x"01",x"23",x"7E",x"FD",x"77",x"02",x"23", -- 0x03E0
    x"7E",x"FD",x"77",x"03",x"F5",x"FD",x"5E",x"00", -- 0x03E8
    x"FD",x"56",x"01",x"FD",x"4E",x"02",x"FD",x"6E", -- 0x03F0
    x"03",x"F1",x"06",x"09",x"CB",x"3D",x"CB",x"19", -- 0x03F8
    x"CB",x"1A",x"CB",x"1B",x"10",x"F6",x"FD",x"21", -- 0x0400
    x"02",x"00",x"FD",x"39",x"FD",x"73",x"00",x"FD", -- 0x0408
    x"72",x"01",x"FD",x"7E",x"00",x"87",x"47",x"0E", -- 0x0410
    x"00",x"11",x"00",x"00",x"21",x"14",x"00",x"39", -- 0x0418
    x"79",x"96",x"78",x"23",x"9E",x"7B",x"23",x"9E", -- 0x0420
    x"7A",x"23",x"9E",x"30",x"08",x"FD",x"34",x"00", -- 0x0428
    x"20",x"03",x"FD",x"34",x"01",x"21",x"3F",x"01", -- 0x0430
    x"4E",x"21",x"02",x"F8",x"71",x"E5",x"CD",x"BB", -- 0x0438
    x"08",x"F1",x"FD",x"21",x"65",x"FC",x"FD",x"75", -- 0x0440
    x"00",x"FD",x"7E",x"00",x"D6",x"12",x"28",x"1D", -- 0x0448
    x"FD",x"7E",x"00",x"D6",x"15",x"28",x"16",x"FD", -- 0x0450
    x"7E",x"00",x"D6",x"16",x"28",x"0F",x"FD",x"7E", -- 0x0458
    x"00",x"D6",x"17",x"28",x"08",x"21",x"E8",x"06", -- 0x0460
    x"E5",x"CD",x"03",x"01",x"F1",x"21",x"02",x"04", -- 0x0468
    x"E5",x"CD",x"2A",x"1E",x"21",x"FF",x"06",x"E3", -- 0x0470
    x"CD",x"B4",x"1F",x"21",x"02",x"06",x"E3",x"CD", -- 0x0478
    x"2A",x"1E",x"21",x"1B",x"07",x"E3",x"CD",x"B4", -- 0x0480
    x"1F",x"F1",x"21",x"3B",x"01",x"46",x"C5",x"33", -- 0x0488
    x"CD",x"F5",x"08",x"33",x"21",x"43",x"01",x"46", -- 0x0490
    x"C5",x"33",x"CD",x"F5",x"08",x"33",x"21",x"65", -- 0x0498
    x"FC",x"36",x"00",x"21",x"3D",x"01",x"46",x"C5", -- 0x04A0
    x"33",x"CD",x"0A",x"09",x"33",x"7D",x"E6",x"01", -- 0x04A8
    x"3D",x"C2",x"38",x"05",x"3E",x"36",x"21",x"65", -- 0x04B0
    x"FC",x"FD",x"21",x"14",x"00",x"FD",x"39",x"86", -- 0x04B8
    x"FD",x"77",x"00",x"3E",x"01",x"CE",x"00",x"FD", -- 0x04C0
    x"23",x"FD",x"77",x"00",x"21",x"14",x"00",x"39", -- 0x04C8
    x"7E",x"23",x"66",x"6F",x"46",x"C5",x"33",x"CD", -- 0x04D0
    x"4B",x"1E",x"33",x"3E",x"08",x"F5",x"33",x"CD", -- 0x04D8
    x"4B",x"1E",x"33",x"FD",x"21",x"65",x"FC",x"FD", -- 0x04E0
    x"7E",x"00",x"3C",x"E6",x"03",x"FD",x"77",x"00", -- 0x04E8
    x"21",x"04",x"00",x"39",x"36",x"88",x"23",x"36", -- 0x04F0
    x"13",x"21",x"14",x"00",x"39",x"FD",x"21",x"04", -- 0x04F8
    x"00",x"FD",x"39",x"FD",x"7E",x"00",x"C6",x"FF", -- 0x0500
    x"77",x"FD",x"7E",x"01",x"CE",x"FF",x"23",x"77", -- 0x0508
    x"21",x"14",x"00",x"39",x"7E",x"FD",x"21",x"04", -- 0x0510
    x"00",x"FD",x"39",x"FD",x"77",x"00",x"21",x"15", -- 0x0518
    x"00",x"39",x"7E",x"FD",x"21",x"04",x"00",x"FD", -- 0x0520
    x"39",x"FD",x"77",x"01",x"21",x"15",x"00",x"39", -- 0x0528
    x"7E",x"2B",x"B6",x"20",x"C4",x"C3",x"A3",x"04", -- 0x0530
    x"21",x"2B",x"07",x"E5",x"CD",x"B4",x"1F",x"21", -- 0x0538
    x"02",x"08",x"E3",x"CD",x"2A",x"1E",x"21",x"30", -- 0x0540
    x"07",x"E3",x"CD",x"B4",x"1F",x"F1",x"AF",x"FD", -- 0x0548
    x"21",x"28",x"FA",x"FD",x"77",x"00",x"FD",x"77", -- 0x0550
    x"01",x"FD",x"77",x"02",x"FD",x"77",x"03",x"21", -- 0x0558
    x"65",x"FC",x"36",x"00",x"21",x"12",x"00",x"39", -- 0x0560
    x"7E",x"FD",x"21",x"14",x"00",x"FD",x"39",x"FD", -- 0x0568
    x"77",x"00",x"21",x"13",x"00",x"39",x"7E",x"FD", -- 0x0570
    x"21",x"14",x"00",x"FD",x"39",x"FD",x"77",x"01", -- 0x0578
    x"01",x"00",x"00",x"21",x"02",x"00",x"39",x"79", -- 0x0580
    x"96",x"78",x"23",x"9E",x"30",x"5A",x"21",x"14", -- 0x0588
    x"00",x"39",x"5E",x"23",x"56",x"C5",x"21",x"02", -- 0x0590
    x"00",x"39",x"4E",x"23",x"46",x"C5",x"D5",x"CD", -- 0x0598
    x"70",x"19",x"F1",x"F1",x"C1",x"03",x"C5",x"21", -- 0x05A0
    x"00",x"60",x"E5",x"CD",x"CB",x"01",x"F1",x"C1", -- 0x05A8
    x"21",x"28",x"FA",x"7E",x"C6",x"00",x"77",x"23", -- 0x05B0
    x"7E",x"CE",x"01",x"77",x"23",x"7E",x"CE",x"00", -- 0x05B8
    x"77",x"23",x"7E",x"CE",x"00",x"77",x"C5",x"21", -- 0x05C0
    x"00",x"61",x"E5",x"CD",x"CB",x"01",x"F1",x"C1", -- 0x05C8
    x"21",x"28",x"FA",x"7E",x"C6",x"00",x"77",x"23", -- 0x05D0
    x"7E",x"CE",x"01",x"77",x"23",x"7E",x"CE",x"00", -- 0x05D8
    x"77",x"23",x"7E",x"CE",x"00",x"77",x"18",x"9B", -- 0x05E0
    x"21",x"2B",x"07",x"E5",x"CD",x"B4",x"1F",x"F1", -- 0x05E8
    x"21",x"3C",x"01",x"46",x"C5",x"33",x"CD",x"F5", -- 0x05F0
    x"08",x"33",x"3E",x"FF",x"D3",x"E7",x"CD",x"05", -- 0x05F8
    x"1E",x"3E",x"04",x"D3",x"FE",x"21",x"0B",x"09", -- 0x0600
    x"E5",x"CD",x"2A",x"1E",x"21",x"40",x"07",x"E3", -- 0x0608
    x"CD",x"B4",x"1F",x"21",x"07",x"0D",x"E3",x"CD", -- 0x0610
    x"2A",x"1E",x"21",x"4B",x"07",x"E3",x"CD",x"B4", -- 0x0618
    x"1F",x"F1",x"18",x"FE",x"21",x"18",x"00",x"39", -- 0x0620
    x"F9",x"C9",x"4D",x"75",x"6C",x"74",x"69",x"63", -- 0x0628
    x"6F",x"72",x"65",x"20",x"32",x"20",x"43",x"4F", -- 0x0630
    x"52",x"45",x"20",x"75",x"70",x"64",x"61",x"74", -- 0x0638
    x"65",x"72",x"00",x"41",x"54",x"54",x"45",x"4E", -- 0x0640
    x"54",x"49",x"4F",x"4E",x"21",x"00",x"54",x"68", -- 0x0648
    x"65",x"20",x"63",x"6F",x"72",x"65",x"20",x"77", -- 0x0650
    x"69",x"6C",x"6C",x"20",x"62",x"65",x"20",x"6F", -- 0x0658
    x"76",x"65",x"72",x"77",x"72",x"69",x"74",x"74", -- 0x0660
    x"65",x"6E",x"00",x"50",x"72",x"65",x"73",x"73", -- 0x0668
    x"20",x"45",x"4E",x"54",x"45",x"52",x"20",x"77", -- 0x0670
    x"68",x"65",x"6E",x"20",x"72",x"65",x"61",x"64", -- 0x0678
    x"79",x"00",x"56",x"20",x"31",x"2E",x"30",x"31", -- 0x0680
    x"00",x"41",x"72",x"65",x"20",x"79",x"6F",x"75", -- 0x0688
    x"20",x"73",x"75",x"72",x"65",x"3F",x"20",x"28", -- 0x0690
    x"59",x"2F",x"4E",x"29",x"00",x"46",x"61",x"69", -- 0x0698
    x"6C",x"20",x"74",x"6F",x"20",x"69",x"6E",x"69", -- 0x06A0
    x"74",x"20",x"74",x"68",x"65",x"20",x"53",x"44", -- 0x06A8
    x"20",x"63",x"61",x"72",x"64",x"00",x"46",x"61", -- 0x06B0
    x"69",x"6C",x"20",x"74",x"6F",x"20",x"6D",x"6F", -- 0x06B8
    x"75",x"6E",x"74",x"20",x"74",x"68",x"65",x"20", -- 0x06C0
    x"53",x"44",x"20",x"63",x"61",x"72",x"64",x"00", -- 0x06C8
    x"46",x"61",x"69",x"6C",x"20",x"74",x"6F",x"20", -- 0x06D0
    x"6F",x"70",x"65",x"6E",x"20",x"55",x"50",x"44", -- 0x06D8
    x"41",x"54",x"45",x"2E",x"43",x"4F",x"52",x"00", -- 0x06E0
    x"46",x"6C",x"61",x"73",x"68",x"20",x"49",x"43", -- 0x06E8
    x"20",x"6E",x"6F",x"74",x"20",x"64",x"65",x"74", -- 0x06F0
    x"65",x"63",x"74",x"65",x"64",x"21",x"00",x"46", -- 0x06F8
    x"6C",x"61",x"73",x"68",x"20",x"49",x"43",x"20", -- 0x0700
    x"64",x"65",x"74",x"65",x"63",x"74",x"65",x"64", -- 0x0708
    x"3A",x"20",x"57",x"32",x"35",x"51",x"36",x"34", -- 0x0710
    x"42",x"56",x"00",x"45",x"72",x"61",x"73",x"69", -- 0x0718
    x"6E",x"67",x"20",x"46",x"6C",x"61",x"73",x"68", -- 0x0720
    x"3A",x"20",x"00",x"20",x"4F",x"4B",x"0A",x"00", -- 0x0728
    x"57",x"72",x"69",x"74",x"69",x"6E",x"67",x"20", -- 0x0730
    x"46",x"6C",x"61",x"73",x"68",x"3A",x"20",x"00", -- 0x0738
    x"55",x"50",x"44",x"41",x"54",x"45",x"20",x"4F", -- 0x0740
    x"4B",x"21",x"00",x"54",x"75",x"72",x"6E",x"20", -- 0x0748
    x"6F",x"66",x"66",x"20",x"74",x"68",x"65",x"20", -- 0x0750
    x"70",x"6F",x"77",x"65",x"72",x"00",x"55",x"50", -- 0x0758
    x"44",x"41",x"54",x"45",x"20",x"20",x"43",x"4F", -- 0x0760
    x"52",x"00",x"3E",x"FF",x"D3",x"E7",x"06",x"0A", -- 0x0768
    x"3E",x"FF",x"D3",x"EB",x"10",x"FA",x"3E",x"FE", -- 0x0770
    x"D3",x"E7",x"06",x"10",x"3E",x"40",x"11",x"00", -- 0x0778
    x"00",x"C5",x"CD",x"52",x"08",x"C1",x"D2",x"92", -- 0x0780
    x"07",x"10",x"F1",x"2E",x"00",x"3E",x"FF",x"D3", -- 0x0788
    x"E7",x"C9",x"3E",x"48",x"11",x"AA",x"01",x"CD", -- 0x0790
    x"5F",x"08",x"21",x"36",x"08",x"38",x"03",x"21", -- 0x0798
    x"44",x"08",x"01",x"78",x"00",x"C5",x"CD",x"B9", -- 0x07A0
    x"07",x"C1",x"D2",x"BA",x"07",x"10",x"F6",x"0D", -- 0x07A8
    x"20",x"F3",x"2E",x"00",x"3E",x"FF",x"D3",x"E7", -- 0x07B0
    x"C9",x"E9",x"3E",x"7A",x"11",x"00",x"00",x"CD", -- 0x07B8
    x"5F",x"08",x"DA",x"B2",x"07",x"78",x"E6",x"40", -- 0x07C0
    x"32",x"2C",x"FA",x"CC",x"DD",x"07",x"3E",x"FF", -- 0x07C8
    x"D3",x"E7",x"3A",x"2C",x"FA",x"2E",x"03",x"FE", -- 0x07D0
    x"40",x"C8",x"2E",x"02",x"C9",x"3E",x"50",x"01", -- 0x07D8
    x"00",x"00",x"11",x"00",x"02",x"C3",x"3D",x"08", -- 0x07E0
    x"FD",x"21",x"00",x"00",x"FD",x"39",x"FD",x"5E", -- 0x07E8
    x"02",x"FD",x"56",x"03",x"FD",x"4E",x"04",x"FD", -- 0x07F0
    x"46",x"05",x"FD",x"6E",x"06",x"FD",x"66",x"07", -- 0x07F8
    x"3E",x"FE",x"D3",x"E7",x"3A",x"2C",x"FA",x"B7", -- 0x0800
    x"CC",x"2A",x"08",x"3E",x"51",x"CD",x"3D",x"08", -- 0x0808
    x"30",x"03",x"2E",x"00",x"C9",x"CD",x"9F",x"08", -- 0x0810
    x"38",x"F8",x"01",x"EB",x"00",x"ED",x"B2",x"ED", -- 0x0818
    x"B2",x"00",x"DB",x"EB",x"00",x"DB",x"EB",x"2E", -- 0x0820
    x"01",x"C9",x"41",x"4A",x"53",x"1E",x"00",x"CB", -- 0x0828
    x"22",x"CB",x"11",x"CB",x"10",x"C9",x"3E",x"41", -- 0x0830
    x"01",x"00",x"00",x"50",x"59",x"CD",x"78",x"08", -- 0x0838
    x"B7",x"C8",x"37",x"C9",x"3E",x"77",x"CD",x"38", -- 0x0840
    x"08",x"3E",x"69",x"01",x"00",x"40",x"51",x"59", -- 0x0848
    x"18",x"EB",x"01",x"00",x"00",x"CD",x"78",x"08", -- 0x0850
    x"47",x"E6",x"FE",x"78",x"20",x"E4",x"C9",x"CD", -- 0x0858
    x"52",x"08",x"D8",x"F5",x"CD",x"AD",x"08",x"67", -- 0x0860
    x"CD",x"AD",x"08",x"6F",x"CD",x"AD",x"08",x"57", -- 0x0868
    x"CD",x"AD",x"08",x"5F",x"44",x"4D",x"F1",x"C9", -- 0x0870
    x"D3",x"EB",x"F5",x"78",x"00",x"D3",x"EB",x"79", -- 0x0878
    x"00",x"D3",x"EB",x"7A",x"00",x"D3",x"EB",x"7B", -- 0x0880
    x"00",x"D3",x"EB",x"F1",x"FE",x"40",x"06",x"95", -- 0x0888
    x"28",x"08",x"FE",x"48",x"06",x"87",x"28",x"02", -- 0x0890
    x"06",x"FF",x"78",x"D3",x"EB",x"18",x"0E",x"06", -- 0x0898
    x"0A",x"C5",x"CD",x"AD",x"08",x"C1",x"FE",x"FE", -- 0x08A0
    x"C8",x"10",x"F6",x"37",x"C9",x"01",x"64",x"00", -- 0x08A8
    x"DB",x"EB",x"FE",x"FF",x"C0",x"10",x"F9",x"0D", -- 0x08B0
    x"20",x"F6",x"C9",x"C1",x"E1",x"E5",x"C5",x"0E", -- 0x08B8
    x"EB",x"3E",x"7F",x"D3",x"E7",x"ED",x"A3",x"ED", -- 0x08C0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"78",x"00", -- 0x08C8
    x"ED",x"78",x"00",x"ED",x"78",x"6F",x"3E",x"FF", -- 0x08D0
    x"D3",x"E7",x"C9",x"3E",x"7F",x"D3",x"E7",x"3E", -- 0x08D8
    x"AB",x"D3",x"EB",x"00",x"D3",x"EB",x"00",x"D3", -- 0x08E0
    x"EB",x"00",x"D3",x"EB",x"00",x"DB",x"EB",x"6F", -- 0x08E8
    x"3E",x"FF",x"D3",x"E7",x"C9",x"FD",x"21",x"00", -- 0x08F0
    x"00",x"FD",x"39",x"FD",x"6E",x"02",x"3E",x"7F", -- 0x08F8
    x"D3",x"E7",x"7D",x"D3",x"EB",x"3E",x"FF",x"D3", -- 0x0900
    x"E7",x"C9",x"21",x"02",x"00",x"39",x"6E",x"0E", -- 0x0908
    x"EB",x"3E",x"7F",x"D3",x"E7",x"7D",x"ED",x"79", -- 0x0910
    x"00",x"ED",x"78",x"00",x"ED",x"68",x"3E",x"FF", -- 0x0918
    x"D3",x"E7",x"C9",x"C1",x"E1",x"E5",x"C5",x"0E", -- 0x0920
    x"EB",x"3E",x"7F",x"D3",x"E7",x"ED",x"A3",x"ED", -- 0x0928
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0930
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0938
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0940
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0948
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0950
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0958
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0960
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0968
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0970
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0978
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0980
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0988
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0990
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0998
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09A0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09A8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09B0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09B8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09C0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09C8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09D0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09D8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09E0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09E8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09F0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x09F8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A00
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A08
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A10
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A18
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A20
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A28
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A30
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A38
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A40
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A48
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A50
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A58
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A60
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A68
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A70
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A78
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A80
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A88
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A90
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0A98
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AA0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AA8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AB0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AB8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AC0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AC8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AD0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AD8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AE0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AE8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AF0
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0AF8
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0B00
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0B08
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0B10
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0B18
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0B20
    x"A3",x"ED",x"A3",x"ED",x"A3",x"ED",x"A3",x"ED", -- 0x0B28
    x"A3",x"ED",x"A3",x"ED",x"A3",x"3E",x"FF",x"D3", -- 0x0B30
    x"E7",x"C9",x"F5",x"F5",x"F5",x"F5",x"FD",x"21", -- 0x0B38
    x"2D",x"FA",x"FD",x"7E",x"01",x"FD",x"B6",x"00", -- 0x0B40
    x"28",x"5C",x"F5",x"21",x"0C",x"00",x"39",x"7E", -- 0x0B48
    x"FD",x"21",x"02",x"00",x"FD",x"39",x"FD",x"77", -- 0x0B50
    x"00",x"21",x"0D",x"00",x"39",x"7E",x"FD",x"21", -- 0x0B58
    x"02",x"00",x"FD",x"39",x"FD",x"77",x"01",x"21", -- 0x0B60
    x"0E",x"00",x"39",x"7E",x"FD",x"21",x"02",x"00", -- 0x0B68
    x"FD",x"39",x"FD",x"77",x"02",x"21",x"0F",x"00", -- 0x0B70
    x"39",x"7E",x"FD",x"21",x"02",x"00",x"FD",x"39", -- 0x0B78
    x"FD",x"77",x"03",x"F1",x"06",x"07",x"FD",x"CB", -- 0x0B80
    x"03",x"3E",x"FD",x"CB",x"02",x"1E",x"FD",x"CB", -- 0x0B88
    x"01",x"1E",x"FD",x"CB",x"00",x"1E",x"10",x"EE", -- 0x0B90
    x"21",x"0A",x"00",x"39",x"5E",x"CB",x"BB",x"16", -- 0x0B98
    x"00",x"01",x"00",x"00",x"18",x"58",x"F5",x"21", -- 0x0BA0
    x"0C",x"00",x"39",x"7E",x"FD",x"21",x"02",x"00", -- 0x0BA8
    x"FD",x"39",x"FD",x"77",x"00",x"21",x"0D",x"00", -- 0x0BB0
    x"39",x"7E",x"FD",x"21",x"02",x"00",x"FD",x"39", -- 0x0BB8
    x"FD",x"77",x"01",x"21",x"0E",x"00",x"39",x"7E", -- 0x0BC0
    x"FD",x"21",x"02",x"00",x"FD",x"39",x"FD",x"77", -- 0x0BC8
    x"02",x"21",x"0F",x"00",x"39",x"7E",x"FD",x"21", -- 0x0BD0
    x"02",x"00",x"FD",x"39",x"FD",x"77",x"03",x"F1", -- 0x0BD8
    x"06",x"08",x"FD",x"CB",x"03",x"3E",x"FD",x"CB", -- 0x0BE0
    x"02",x"1E",x"FD",x"CB",x"01",x"1E",x"FD",x"CB", -- 0x0BE8
    x"00",x"1E",x"10",x"EE",x"21",x"0A",x"00",x"39", -- 0x0BF0
    x"5E",x"16",x"00",x"01",x"00",x"00",x"21",x"00", -- 0x0BF8
    x"00",x"39",x"7E",x"FD",x"21",x"57",x"FC",x"FD", -- 0x0C00
    x"96",x"00",x"20",x"2A",x"21",x"01",x"00",x"39", -- 0x0C08
    x"7E",x"FD",x"21",x"57",x"FC",x"FD",x"96",x"01", -- 0x0C10
    x"20",x"1C",x"21",x"02",x"00",x"39",x"7E",x"FD", -- 0x0C18
    x"21",x"57",x"FC",x"FD",x"96",x"02",x"20",x"0E", -- 0x0C20
    x"21",x"03",x"00",x"39",x"7E",x"FD",x"21",x"57", -- 0x0C28
    x"FC",x"FD",x"96",x"03",x"28",x"6A",x"21",x"00", -- 0x0C30
    x"00",x"39",x"D5",x"FD",x"21",x"06",x"00",x"FD", -- 0x0C38
    x"39",x"FD",x"E5",x"D1",x"FD",x"21",x"2F",x"FA", -- 0x0C40
    x"FD",x"7E",x"00",x"86",x"12",x"FD",x"7E",x"01", -- 0x0C48
    x"23",x"8E",x"13",x"12",x"FD",x"7E",x"02",x"23", -- 0x0C50
    x"8E",x"13",x"12",x"FD",x"7E",x"03",x"23",x"8E", -- 0x0C58
    x"13",x"12",x"D1",x"C5",x"D5",x"21",x"55",x"FA", -- 0x0C60
    x"E5",x"FD",x"21",x"0A",x"00",x"FD",x"39",x"FD", -- 0x0C68
    x"6E",x"02",x"FD",x"66",x"03",x"E5",x"FD",x"6E", -- 0x0C70
    x"00",x"FD",x"66",x"01",x"E5",x"CD",x"E8",x"07", -- 0x0C78
    x"F1",x"F1",x"F1",x"D1",x"C1",x"7D",x"B7",x"20", -- 0x0C80
    x"07",x"21",x"00",x"00",x"5D",x"54",x"18",x"4D", -- 0x0C88
    x"D5",x"C5",x"11",x"57",x"FC",x"21",x"04",x"00", -- 0x0C90
    x"39",x"01",x"04",x"00",x"ED",x"B0",x"C1",x"D1", -- 0x0C98
    x"FD",x"21",x"2D",x"FA",x"FD",x"7E",x"01",x"FD", -- 0x0CA0
    x"B6",x"00",x"28",x"1D",x"21",x"55",x"FA",x"3E", -- 0x0CA8
    x"02",x"CB",x"23",x"CB",x"12",x"CB",x"11",x"CB", -- 0x0CB0
    x"10",x"3D",x"20",x"F5",x"19",x"4E",x"23",x"46", -- 0x0CB8
    x"23",x"5E",x"23",x"7E",x"E6",x"0F",x"57",x"18", -- 0x0CC0
    x"12",x"21",x"55",x"FA",x"CB",x"23",x"CB",x"12", -- 0x0CC8
    x"CB",x"11",x"CB",x"10",x"19",x"4E",x"23",x"46", -- 0x0CD0
    x"11",x"00",x"00",x"69",x"60",x"F1",x"F1",x"F1", -- 0x0CD8
    x"F1",x"C9",x"F5",x"F5",x"21",x"06",x"00",x"39", -- 0x0CE0
    x"4E",x"23",x"46",x"21",x"08",x"00",x"39",x"7E", -- 0x0CE8
    x"FD",x"21",x"02",x"00",x"FD",x"39",x"FD",x"77", -- 0x0CF0
    x"00",x"21",x"09",x"00",x"39",x"7E",x"FD",x"21", -- 0x0CF8
    x"02",x"00",x"FD",x"39",x"FD",x"77",x"01",x"11", -- 0x0D00
    x"00",x"00",x"21",x"0A",x"00",x"39",x"7B",x"96", -- 0x0D08
    x"7A",x"23",x"9E",x"E2",x"18",x"0D",x"EE",x"80", -- 0x0D10
    x"F2",x"58",x"0D",x"0A",x"33",x"F5",x"33",x"03", -- 0x0D18
    x"21",x"02",x"00",x"39",x"7E",x"23",x"66",x"6F", -- 0x0D20
    x"7E",x"FD",x"21",x"01",x"00",x"FD",x"39",x"FD", -- 0x0D28
    x"77",x"00",x"FD",x"21",x"02",x"00",x"FD",x"39", -- 0x0D30
    x"FD",x"34",x"00",x"20",x"03",x"FD",x"34",x"01", -- 0x0D38
    x"21",x"00",x"00",x"39",x"7E",x"FD",x"21",x"01", -- 0x0D40
    x"00",x"FD",x"39",x"FD",x"96",x"00",x"28",x"05", -- 0x0D48
    x"21",x"01",x"00",x"18",x"06",x"13",x"18",x"B2", -- 0x0D50
    x"21",x"00",x"00",x"F1",x"F1",x"C9",x"21",x"F5", -- 0x0D58
    x"FF",x"39",x"F9",x"FD",x"21",x"57",x"FC",x"FD", -- 0x0D60
    x"36",x"00",x"FF",x"FD",x"36",x"01",x"FF",x"FD", -- 0x0D68
    x"36",x"02",x"FF",x"FD",x"36",x"03",x"FF",x"21", -- 0x0D70
    x"00",x"00",x"22",x"2D",x"FA",x"21",x"55",x"FA", -- 0x0D78
    x"E5",x"21",x"00",x"00",x"E5",x"21",x"00",x"00", -- 0x0D80
    x"E5",x"CD",x"E8",x"07",x"F1",x"F1",x"F1",x"FD", -- 0x0D88
    x"21",x"0A",x"00",x"FD",x"39",x"FD",x"75",x"00", -- 0x0D90
    x"21",x"0A",x"00",x"39",x"7E",x"B7",x"20",x"04", -- 0x0D98
    x"6F",x"C3",x"A3",x"15",x"AF",x"FD",x"21",x"06", -- 0x0DA0
    x"00",x"FD",x"39",x"FD",x"77",x"00",x"FD",x"77", -- 0x0DA8
    x"01",x"FD",x"77",x"02",x"FD",x"77",x"03",x"21", -- 0x0DB0
    x"01",x"00",x"22",x"55",x"FC",x"2E",x"08",x"E5", -- 0x0DB8
    x"21",x"AC",x"15",x"E5",x"21",x"8B",x"FA",x"E5", -- 0x0DC0
    x"CD",x"E2",x"0C",x"F1",x"F1",x"F1",x"7C",x"B5", -- 0x0DC8
    x"20",x"06",x"21",x"00",x"00",x"22",x"55",x"FC", -- 0x0DD0
    x"21",x"08",x"00",x"E5",x"21",x"B5",x"15",x"E5", -- 0x0DD8
    x"21",x"A7",x"FA",x"E5",x"CD",x"E2",x"0C",x"F1", -- 0x0DE0
    x"F1",x"F1",x"7C",x"B5",x"20",x"06",x"21",x"00", -- 0x0DE8
    x"00",x"22",x"55",x"FC",x"FD",x"21",x"55",x"FC", -- 0x0DF0
    x"FD",x"7E",x"01",x"FD",x"B6",x"00",x"CA",x"7E", -- 0x0DF8
    x"0E",x"01",x"55",x"FA",x"33",x"33",x"C5",x"E1", -- 0x0E00
    x"E5",x"11",x"C6",x"01",x"19",x"4E",x"23",x"46", -- 0x0E08
    x"23",x"5E",x"23",x"56",x"FD",x"21",x"06",x"00", -- 0x0E10
    x"FD",x"39",x"FD",x"71",x"00",x"FD",x"70",x"01", -- 0x0E18
    x"FD",x"73",x"02",x"FD",x"72",x"03",x"E1",x"E5", -- 0x0E20
    x"C5",x"01",x"FE",x"01",x"09",x"C1",x"7E",x"23", -- 0x0E28
    x"66",x"6F",x"D6",x"AA",x"20",x"13",x"7C",x"D6", -- 0x0E30
    x"55",x"20",x"0E",x"FD",x"71",x"00",x"FD",x"70", -- 0x0E38
    x"01",x"FD",x"73",x"02",x"FD",x"72",x"03",x"18", -- 0x0E40
    x"0F",x"7D",x"D6",x"55",x"20",x"05",x"7C",x"D6", -- 0x0E48
    x"AA",x"28",x"05",x"2E",x"00",x"C3",x"A3",x"15", -- 0x0E50
    x"21",x"55",x"FA",x"E5",x"FD",x"21",x"08",x"00", -- 0x0E58
    x"FD",x"39",x"FD",x"6E",x"02",x"FD",x"66",x"03", -- 0x0E60
    x"E5",x"FD",x"6E",x"00",x"FD",x"66",x"01",x"E5", -- 0x0E68
    x"CD",x"E8",x"07",x"F1",x"F1",x"F1",x"7D",x"B7", -- 0x0E70
    x"20",x"04",x"6F",x"C3",x"A3",x"15",x"21",x"08", -- 0x0E78
    x"00",x"E5",x"21",x"B5",x"15",x"E5",x"21",x"A7", -- 0x0E80
    x"FA",x"E5",x"CD",x"E2",x"0C",x"F1",x"F1",x"F1", -- 0x0E88
    x"7C",x"B5",x"20",x"08",x"21",x"01",x"00",x"22", -- 0x0E90
    x"2D",x"FA",x"18",x"1B",x"21",x"08",x"00",x"E5", -- 0x0E98
    x"21",x"AC",x"15",x"E5",x"21",x"8B",x"FA",x"E5", -- 0x0EA0
    x"CD",x"E2",x"0C",x"F1",x"F1",x"F1",x"7C",x"B5", -- 0x0EA8
    x"28",x"05",x"2E",x"00",x"C3",x"A3",x"15",x"3A", -- 0x0EB0
    x"53",x"FC",x"D6",x"55",x"20",x"07",x"3A",x"54", -- 0x0EB8
    x"FC",x"D6",x"AA",x"28",x"05",x"2E",x"00",x"C3", -- 0x0EC0
    x"A3",x"15",x"21",x"55",x"FA",x"4E",x"79",x"FE", -- 0x0EC8
    x"E9",x"28",x"09",x"D6",x"EB",x"28",x"05",x"2E", -- 0x0ED0
    x"00",x"C3",x"A3",x"15",x"3A",x"60",x"FA",x"B7", -- 0x0ED8
    x"20",x"07",x"3A",x"61",x"FA",x"D6",x"02",x"28", -- 0x0EE0
    x"05",x"2E",x"00",x"C3",x"A3",x"15",x"3A",x"62", -- 0x0EE8
    x"FA",x"FD",x"21",x"45",x"FA",x"FD",x"77",x"00", -- 0x0EF0
    x"FD",x"36",x"01",x"00",x"FD",x"36",x"02",x"00", -- 0x0EF8
    x"FD",x"36",x"03",x"00",x"21",x"49",x"FA",x"FD", -- 0x0F00
    x"7E",x"00",x"C6",x"FF",x"77",x"FD",x"7E",x"01", -- 0x0F08
    x"CE",x"FF",x"23",x"77",x"FD",x"7E",x"02",x"CE", -- 0x0F10
    x"FF",x"23",x"77",x"FD",x"7E",x"03",x"CE",x"FF", -- 0x0F18
    x"23",x"77",x"3A",x"63",x"FA",x"FD",x"21",x"0A", -- 0x0F20
    x"00",x"FD",x"39",x"FD",x"77",x"00",x"FD",x"7E", -- 0x0F28
    x"00",x"FD",x"21",x"02",x"00",x"FD",x"39",x"FD", -- 0x0F30
    x"77",x"00",x"FD",x"36",x"01",x"00",x"FD",x"36", -- 0x0F38
    x"02",x"00",x"FD",x"36",x"03",x"00",x"21",x"02", -- 0x0F40
    x"00",x"39",x"FD",x"21",x"06",x"00",x"FD",x"39", -- 0x0F48
    x"FD",x"7E",x"00",x"86",x"77",x"FD",x"7E",x"01", -- 0x0F50
    x"23",x"8E",x"77",x"FD",x"7E",x"02",x"23",x"8E", -- 0x0F58
    x"77",x"FD",x"7E",x"03",x"23",x"8E",x"77",x"3A", -- 0x0F60
    x"64",x"FA",x"FD",x"77",x"00",x"FD",x"7E",x"00", -- 0x0F68
    x"FD",x"77",x"00",x"FD",x"36",x"01",x"00",x"FD", -- 0x0F70
    x"7E",x"00",x"FD",x"77",x"01",x"FD",x"36",x"00", -- 0x0F78
    x"00",x"FD",x"7E",x"00",x"FD",x"77",x"00",x"FD", -- 0x0F80
    x"7E",x"01",x"FD",x"77",x"01",x"FD",x"7E",x"01", -- 0x0F88
    x"17",x"9F",x"FD",x"77",x"02",x"FD",x"77",x"03", -- 0x0F90
    x"21",x"06",x"00",x"39",x"D5",x"11",x"2F",x"FA", -- 0x0F98
    x"FD",x"21",x"04",x"00",x"FD",x"39",x"FD",x"7E", -- 0x0FA0
    x"00",x"86",x"12",x"FD",x"7E",x"01",x"23",x"8E", -- 0x0FA8
    x"13",x"12",x"FD",x"7E",x"02",x"23",x"8E",x"13", -- 0x0FB0
    x"12",x"FD",x"7E",x"03",x"23",x"8E",x"13",x"12", -- 0x0FB8
    x"D1",x"3A",x"65",x"FA",x"FD",x"21",x"43",x"FA", -- 0x0FC0
    x"FD",x"77",x"00",x"FD",x"36",x"01",x"00",x"FD", -- 0x0FC8
    x"21",x"2D",x"FA",x"FD",x"7E",x"01",x"FD",x"B6", -- 0x0FD0
    x"00",x"CA",x"8B",x"13",x"21",x"08",x"00",x"E5", -- 0x0FD8
    x"21",x"B5",x"15",x"E5",x"21",x"A7",x"FA",x"E5", -- 0x0FE0
    x"CD",x"E2",x"0C",x"F1",x"F1",x"F1",x"7C",x"B5", -- 0x0FE8
    x"28",x"05",x"2E",x"00",x"C3",x"A3",x"15",x"F5", -- 0x0FF0
    x"3A",x"45",x"FA",x"FD",x"21",x"4D",x"FA",x"FD", -- 0x0FF8
    x"77",x"00",x"3A",x"46",x"FA",x"FD",x"21",x"4D", -- 0x1000
    x"FA",x"FD",x"77",x"01",x"3A",x"47",x"FA",x"FD", -- 0x1008
    x"21",x"4D",x"FA",x"FD",x"77",x"02",x"3A",x"48", -- 0x1010
    x"FA",x"FD",x"21",x"4D",x"FA",x"FD",x"77",x"03", -- 0x1018
    x"F1",x"06",x"04",x"FD",x"CB",x"00",x"26",x"FD", -- 0x1020
    x"CB",x"01",x"16",x"FD",x"CB",x"02",x"16",x"FD", -- 0x1028
    x"CB",x"03",x"16",x"10",x"EE",x"11",x"3F",x"FA", -- 0x1030
    x"21",x"45",x"FA",x"01",x"04",x"00",x"ED",x"B0", -- 0x1038
    x"3A",x"79",x"FA",x"FD",x"21",x"02",x"00",x"FD", -- 0x1040
    x"39",x"FD",x"77",x"00",x"3A",x"7A",x"FA",x"FD", -- 0x1048
    x"21",x"06",x"00",x"FD",x"39",x"FD",x"77",x"00", -- 0x1050
    x"FD",x"7E",x"00",x"FD",x"77",x"00",x"FD",x"36", -- 0x1058
    x"01",x"00",x"FD",x"36",x"02",x"00",x"FD",x"36", -- 0x1060
    x"03",x"00",x"F5",x"F1",x"06",x"08",x"FD",x"CB", -- 0x1068
    x"00",x"26",x"FD",x"CB",x"01",x"16",x"FD",x"CB", -- 0x1070
    x"02",x"16",x"FD",x"CB",x"03",x"16",x"10",x"EE", -- 0x1078
    x"FD",x"21",x"02",x"00",x"FD",x"39",x"FD",x"7E", -- 0x1080
    x"00",x"FD",x"77",x"00",x"FD",x"36",x"01",x"00", -- 0x1088
    x"FD",x"36",x"02",x"00",x"FD",x"36",x"03",x"00", -- 0x1090
    x"21",x"06",x"00",x"39",x"D5",x"FD",x"E5",x"D1", -- 0x1098
    x"1A",x"86",x"12",x"13",x"1A",x"23",x"8E",x"12", -- 0x10A0
    x"13",x"1A",x"23",x"8E",x"12",x"13",x"1A",x"23", -- 0x10A8
    x"8E",x"12",x"D1",x"3A",x"7B",x"FA",x"FD",x"21", -- 0x10B0
    x"06",x"00",x"FD",x"39",x"FD",x"77",x"00",x"FD", -- 0x10B8
    x"7E",x"00",x"FD",x"77",x"00",x"FD",x"36",x"01", -- 0x10C0
    x"00",x"FD",x"36",x"02",x"00",x"FD",x"36",x"03", -- 0x10C8
    x"00",x"F5",x"F1",x"06",x"10",x"FD",x"CB",x"00", -- 0x10D0
    x"26",x"FD",x"CB",x"01",x"16",x"FD",x"CB",x"02", -- 0x10D8
    x"16",x"FD",x"CB",x"03",x"16",x"10",x"EE",x"21", -- 0x10E0
    x"06",x"00",x"39",x"D5",x"FD",x"21",x"04",x"00", -- 0x10E8
    x"FD",x"39",x"FD",x"E5",x"D1",x"1A",x"86",x"12", -- 0x10F0
    x"13",x"1A",x"23",x"8E",x"12",x"13",x"1A",x"23", -- 0x10F8
    x"8E",x"12",x"13",x"1A",x"23",x"8E",x"12",x"D1", -- 0x1100
    x"3A",x"7C",x"FA",x"FD",x"21",x"06",x"00",x"FD", -- 0x1108
    x"39",x"FD",x"77",x"00",x"FD",x"7E",x"00",x"FD", -- 0x1110
    x"77",x"00",x"FD",x"36",x"01",x"00",x"FD",x"36", -- 0x1118
    x"02",x"00",x"FD",x"36",x"03",x"00",x"F5",x"F1", -- 0x1120
    x"06",x"18",x"FD",x"CB",x"00",x"26",x"FD",x"CB", -- 0x1128
    x"01",x"16",x"FD",x"CB",x"02",x"16",x"FD",x"CB", -- 0x1130
    x"03",x"16",x"10",x"EE",x"21",x"06",x"00",x"39", -- 0x1138
    x"D5",x"11",x"51",x"FA",x"FD",x"21",x"04",x"00", -- 0x1140
    x"FD",x"39",x"FD",x"7E",x"00",x"86",x"12",x"FD", -- 0x1148
    x"7E",x"01",x"23",x"8E",x"13",x"12",x"FD",x"7E", -- 0x1150
    x"02",x"23",x"8E",x"13",x"12",x"FD",x"7E",x"03", -- 0x1158
    x"23",x"8E",x"13",x"12",x"D1",x"3A",x"43",x"FA", -- 0x1160
    x"FD",x"21",x"02",x"00",x"FD",x"39",x"FD",x"77", -- 0x1168
    x"00",x"3A",x"44",x"FA",x"FD",x"21",x"02",x"00", -- 0x1170
    x"FD",x"39",x"FD",x"77",x"01",x"FD",x"36",x"02", -- 0x1178
    x"00",x"FD",x"36",x"03",x"00",x"2A",x"53",x"FA", -- 0x1180
    x"E5",x"2A",x"51",x"FA",x"E5",x"FD",x"6E",x"02", -- 0x1188
    x"FD",x"66",x"03",x"E5",x"FD",x"6E",x"00",x"FD", -- 0x1190
    x"66",x"01",x"E5",x"CD",x"7B",x"20",x"F1",x"F1", -- 0x1198
    x"F1",x"F1",x"FD",x"21",x"02",x"00",x"FD",x"39", -- 0x11A0
    x"FD",x"72",x"03",x"FD",x"73",x"02",x"FD",x"74", -- 0x11A8
    x"01",x"FD",x"75",x"00",x"21",x"02",x"00",x"39", -- 0x11B0
    x"D5",x"11",x"33",x"FA",x"FD",x"21",x"2F",x"FA", -- 0x11B8
    x"FD",x"7E",x"00",x"86",x"12",x"FD",x"7E",x"01", -- 0x11C0
    x"23",x"8E",x"13",x"12",x"FD",x"7E",x"02",x"23", -- 0x11C8
    x"8E",x"13",x"12",x"FD",x"7E",x"03",x"23",x"8E", -- 0x11D0
    x"13",x"12",x"D1",x"3A",x"81",x"FA",x"FD",x"21", -- 0x11D8
    x"02",x"00",x"FD",x"39",x"FD",x"77",x"00",x"3A", -- 0x11E0
    x"82",x"FA",x"FD",x"21",x"06",x"00",x"FD",x"39", -- 0x11E8
    x"FD",x"77",x"00",x"FD",x"7E",x"00",x"FD",x"77", -- 0x11F0
    x"00",x"FD",x"36",x"01",x"00",x"FD",x"36",x"02", -- 0x11F8
    x"00",x"FD",x"36",x"03",x"00",x"F5",x"F1",x"06", -- 0x1200
    x"08",x"FD",x"CB",x"00",x"26",x"FD",x"CB",x"01", -- 0x1208
    x"16",x"FD",x"CB",x"02",x"16",x"FD",x"CB",x"03", -- 0x1210
    x"16",x"10",x"EE",x"FD",x"21",x"02",x"00",x"FD", -- 0x1218
    x"39",x"FD",x"7E",x"00",x"FD",x"77",x"00",x"FD", -- 0x1220
    x"36",x"01",x"00",x"FD",x"36",x"02",x"00",x"FD", -- 0x1228
    x"36",x"03",x"00",x"21",x"06",x"00",x"39",x"D5", -- 0x1230
    x"FD",x"E5",x"D1",x"1A",x"86",x"12",x"13",x"1A", -- 0x1238
    x"23",x"8E",x"12",x"13",x"1A",x"23",x"8E",x"12", -- 0x1240
    x"13",x"1A",x"23",x"8E",x"12",x"D1",x"3A",x"83", -- 0x1248
    x"FA",x"FD",x"21",x"06",x"00",x"FD",x"39",x"FD", -- 0x1250
    x"77",x"00",x"FD",x"7E",x"00",x"FD",x"77",x"00", -- 0x1258
    x"FD",x"36",x"01",x"00",x"FD",x"36",x"02",x"00", -- 0x1260
    x"FD",x"36",x"03",x"00",x"F5",x"F1",x"06",x"10", -- 0x1268
    x"FD",x"CB",x"00",x"26",x"FD",x"CB",x"01",x"16", -- 0x1270
    x"FD",x"CB",x"02",x"16",x"FD",x"CB",x"03",x"16", -- 0x1278
    x"10",x"EE",x"21",x"06",x"00",x"39",x"D5",x"FD", -- 0x1280
    x"21",x"04",x"00",x"FD",x"39",x"FD",x"E5",x"D1", -- 0x1288
    x"1A",x"86",x"12",x"13",x"1A",x"23",x"8E",x"12", -- 0x1290
    x"13",x"1A",x"23",x"8E",x"12",x"13",x"1A",x"23", -- 0x1298
    x"8E",x"12",x"D1",x"3A",x"84",x"FA",x"FD",x"21", -- 0x12A0
    x"06",x"00",x"FD",x"39",x"FD",x"77",x"00",x"FD", -- 0x12A8
    x"7E",x"00",x"E6",x"0F",x"FD",x"77",x"00",x"FD", -- 0x12B0
    x"7E",x"00",x"FD",x"77",x"00",x"FD",x"36",x"01", -- 0x12B8
    x"00",x"FD",x"36",x"02",x"00",x"FD",x"36",x"03", -- 0x12C0
    x"00",x"F5",x"F1",x"06",x"18",x"FD",x"CB",x"00", -- 0x12C8
    x"26",x"FD",x"CB",x"01",x"16",x"FD",x"CB",x"02", -- 0x12D0
    x"16",x"FD",x"CB",x"03",x"16",x"10",x"EE",x"21", -- 0x12D8
    x"06",x"00",x"39",x"D5",x"11",x"37",x"FA",x"FD", -- 0x12E0
    x"21",x"04",x"00",x"FD",x"39",x"FD",x"7E",x"00", -- 0x12E8
    x"86",x"12",x"FD",x"7E",x"01",x"23",x"8E",x"13", -- 0x12F0
    x"12",x"FD",x"7E",x"02",x"23",x"8E",x"13",x"12", -- 0x12F8
    x"FD",x"7E",x"03",x"23",x"8E",x"13",x"12",x"D1", -- 0x1300
    x"21",x"02",x"00",x"39",x"FD",x"21",x"37",x"FA", -- 0x1308
    x"FD",x"7E",x"00",x"C6",x"FE",x"77",x"FD",x"7E", -- 0x1310
    x"01",x"CE",x"FF",x"23",x"77",x"FD",x"7E",x"02", -- 0x1318
    x"CE",x"FF",x"23",x"77",x"FD",x"7E",x"03",x"CE", -- 0x1320
    x"FF",x"23",x"77",x"2A",x"47",x"FA",x"E5",x"2A", -- 0x1328
    x"45",x"FA",x"E5",x"FD",x"21",x"06",x"00",x"FD", -- 0x1330
    x"39",x"FD",x"6E",x"02",x"FD",x"66",x"03",x"E5", -- 0x1338
    x"FD",x"6E",x"00",x"FD",x"66",x"01",x"E5",x"CD", -- 0x1340
    x"7B",x"20",x"F1",x"F1",x"F1",x"F1",x"FD",x"21", -- 0x1348
    x"02",x"00",x"FD",x"39",x"FD",x"72",x"03",x"FD", -- 0x1350
    x"73",x"02",x"FD",x"74",x"01",x"FD",x"75",x"00", -- 0x1358
    x"21",x"33",x"FA",x"D5",x"11",x"3B",x"FA",x"FD", -- 0x1360
    x"21",x"04",x"00",x"FD",x"39",x"FD",x"7E",x"00", -- 0x1368
    x"86",x"12",x"FD",x"7E",x"01",x"23",x"8E",x"13", -- 0x1370
    x"12",x"FD",x"7E",x"02",x"23",x"8E",x"13",x"12", -- 0x1378
    x"FD",x"7E",x"03",x"23",x"8E",x"13",x"12",x"D1", -- 0x1380
    x"C3",x"A1",x"15",x"3A",x"66",x"FA",x"FD",x"21", -- 0x1388
    x"02",x"00",x"FD",x"39",x"FD",x"77",x"00",x"FD", -- 0x1390
    x"36",x"01",x"00",x"3A",x"67",x"FA",x"FD",x"21", -- 0x1398
    x"06",x"00",x"FD",x"39",x"FD",x"77",x"00",x"FD", -- 0x13A0
    x"7E",x"00",x"FD",x"77",x"00",x"FD",x"36",x"01", -- 0x13A8
    x"00",x"FD",x"7E",x"00",x"FD",x"77",x"01",x"FD", -- 0x13B0
    x"36",x"00",x"00",x"21",x"06",x"00",x"39",x"D5", -- 0x13B8
    x"FD",x"21",x"04",x"00",x"FD",x"39",x"FD",x"E5", -- 0x13C0
    x"D1",x"FD",x"7E",x"00",x"86",x"12",x"FD",x"7E", -- 0x13C8
    x"01",x"23",x"8E",x"13",x"12",x"D1",x"FD",x"7E", -- 0x13D0
    x"00",x"32",x"4D",x"FA",x"21",x"03",x"00",x"39", -- 0x13D8
    x"7E",x"32",x"4E",x"FA",x"21",x"03",x"00",x"39", -- 0x13E0
    x"7E",x"17",x"9F",x"FD",x"21",x"4D",x"FA",x"FD", -- 0x13E8
    x"77",x"02",x"FD",x"77",x"03",x"F5",x"FD",x"7E", -- 0x13F0
    x"00",x"FD",x"21",x"04",x"00",x"FD",x"39",x"FD", -- 0x13F8
    x"77",x"00",x"3A",x"4E",x"FA",x"FD",x"21",x"04", -- 0x1400
    x"00",x"FD",x"39",x"FD",x"77",x"01",x"3A",x"4F", -- 0x1408
    x"FA",x"FD",x"21",x"04",x"00",x"FD",x"39",x"FD", -- 0x1410
    x"77",x"02",x"3A",x"50",x"FA",x"FD",x"21",x"04", -- 0x1418
    x"00",x"FD",x"39",x"FD",x"77",x"03",x"F1",x"06", -- 0x1420
    x"05",x"FD",x"CB",x"00",x"26",x"FD",x"CB",x"01", -- 0x1428
    x"16",x"FD",x"CB",x"02",x"16",x"FD",x"CB",x"03", -- 0x1430
    x"16",x"10",x"EE",x"21",x"02",x"00",x"39",x"7E", -- 0x1438
    x"C6",x"FF",x"77",x"23",x"7E",x"CE",x"01",x"77", -- 0x1440
    x"23",x"7E",x"CE",x"00",x"77",x"23",x"7E",x"CE", -- 0x1448
    x"00",x"77",x"F5",x"FD",x"7E",x"00",x"32",x"3F", -- 0x1450
    x"FA",x"21",x"05",x"00",x"39",x"7E",x"32",x"40", -- 0x1458
    x"FA",x"21",x"06",x"00",x"39",x"7E",x"32",x"41", -- 0x1460
    x"FA",x"21",x"07",x"00",x"39",x"7E",x"FD",x"21", -- 0x1468
    x"3F",x"FA",x"FD",x"77",x"03",x"F1",x"06",x"09", -- 0x1470
    x"FD",x"CB",x"03",x"3E",x"FD",x"CB",x"02",x"1E", -- 0x1478
    x"FD",x"CB",x"01",x"1E",x"FD",x"CB",x"00",x"1E", -- 0x1480
    x"10",x"EE",x"3A",x"6B",x"FA",x"FD",x"21",x"02", -- 0x1488
    x"00",x"FD",x"39",x"FD",x"77",x"00",x"FD",x"36", -- 0x1490
    x"01",x"00",x"3A",x"6C",x"FA",x"FD",x"21",x"06", -- 0x1498
    x"00",x"FD",x"39",x"FD",x"77",x"00",x"FD",x"7E", -- 0x14A0
    x"00",x"FD",x"77",x"00",x"FD",x"36",x"01",x"00", -- 0x14A8
    x"FD",x"7E",x"00",x"FD",x"77",x"01",x"FD",x"36", -- 0x14B0
    x"00",x"00",x"21",x"06",x"00",x"39",x"D5",x"FD", -- 0x14B8
    x"21",x"04",x"00",x"FD",x"39",x"FD",x"E5",x"D1", -- 0x14C0
    x"FD",x"7E",x"00",x"86",x"12",x"FD",x"7E",x"01", -- 0x14C8
    x"23",x"8E",x"13",x"12",x"D1",x"FD",x"7E",x"00", -- 0x14D0
    x"32",x"51",x"FA",x"21",x"03",x"00",x"39",x"7E", -- 0x14D8
    x"32",x"52",x"FA",x"21",x"03",x"00",x"39",x"7E", -- 0x14E0
    x"17",x"9F",x"FD",x"21",x"51",x"FA",x"FD",x"77", -- 0x14E8
    x"02",x"FD",x"77",x"03",x"3A",x"43",x"FA",x"FD", -- 0x14F0
    x"21",x"02",x"00",x"FD",x"39",x"FD",x"77",x"00", -- 0x14F8
    x"3A",x"44",x"FA",x"FD",x"21",x"02",x"00",x"FD", -- 0x1500
    x"39",x"FD",x"77",x"01",x"FD",x"36",x"02",x"00", -- 0x1508
    x"FD",x"36",x"03",x"00",x"2A",x"53",x"FA",x"E5", -- 0x1510
    x"2A",x"51",x"FA",x"E5",x"FD",x"6E",x"02",x"FD", -- 0x1518
    x"66",x"03",x"E5",x"FD",x"6E",x"00",x"FD",x"66", -- 0x1520
    x"01",x"E5",x"CD",x"7B",x"20",x"F1",x"F1",x"F1", -- 0x1528
    x"F1",x"FD",x"21",x"02",x"00",x"FD",x"39",x"FD", -- 0x1530
    x"72",x"03",x"FD",x"73",x"02",x"FD",x"74",x"01", -- 0x1538
    x"FD",x"75",x"00",x"21",x"02",x"00",x"39",x"D5", -- 0x1540
    x"11",x"3B",x"FA",x"FD",x"21",x"2F",x"FA",x"FD", -- 0x1548
    x"7E",x"00",x"86",x"12",x"FD",x"7E",x"01",x"23", -- 0x1550
    x"8E",x"13",x"12",x"FD",x"7E",x"02",x"23",x"8E", -- 0x1558
    x"13",x"12",x"FD",x"7E",x"03",x"23",x"8E",x"13", -- 0x1560
    x"12",x"D1",x"AF",x"FD",x"21",x"37",x"FA",x"FD", -- 0x1568
    x"77",x"00",x"FD",x"77",x"01",x"FD",x"77",x"02", -- 0x1570
    x"FD",x"77",x"03",x"21",x"3F",x"FA",x"D5",x"11", -- 0x1578
    x"33",x"FA",x"FD",x"21",x"3B",x"FA",x"FD",x"7E", -- 0x1580
    x"00",x"86",x"12",x"FD",x"7E",x"01",x"23",x"8E", -- 0x1588
    x"13",x"12",x"FD",x"7E",x"02",x"23",x"8E",x"13", -- 0x1590
    x"12",x"FD",x"7E",x"03",x"23",x"8E",x"13",x"12", -- 0x1598
    x"D1",x"2E",x"01",x"FD",x"21",x"0B",x"00",x"FD", -- 0x15A0
    x"39",x"FD",x"F9",x"C9",x"46",x"41",x"54",x"31", -- 0x15A8
    x"36",x"20",x"20",x"20",x"00",x"46",x"41",x"54", -- 0x15B0
    x"33",x"32",x"20",x"20",x"20",x"00",x"21",x"E0", -- 0x15B8
    x"FF",x"39",x"F9",x"21",x"0C",x"00",x"39",x"36", -- 0x15C0
    x"00",x"23",x"36",x"00",x"FD",x"21",x"57",x"FC", -- 0x15C8
    x"FD",x"36",x"00",x"FF",x"FD",x"36",x"01",x"FF", -- 0x15D0
    x"FD",x"36",x"02",x"FF",x"FD",x"36",x"03",x"FF", -- 0x15D8
    x"21",x"08",x"00",x"39",x"EB",x"21",x"37",x"FA", -- 0x15E0
    x"01",x"04",x"00",x"ED",x"B0",x"21",x"0E",x"00", -- 0x15E8
    x"39",x"EB",x"21",x"3B",x"FA",x"01",x"04",x"00", -- 0x15F0
    x"ED",x"B0",x"FD",x"21",x"2D",x"FA",x"FD",x"7E", -- 0x15F8
    x"01",x"FD",x"B6",x"00",x"28",x"1E",x"F5",x"FD", -- 0x1600
    x"21",x"45",x"FA",x"FD",x"5E",x"00",x"FD",x"56", -- 0x1608
    x"01",x"FD",x"6E",x"02",x"FD",x"66",x"03",x"F1", -- 0x1610
    x"06",x"04",x"CB",x"23",x"CB",x"12",x"ED",x"6A", -- 0x1618
    x"10",x"F8",x"18",x"1C",x"F5",x"FD",x"21",x"3F", -- 0x1620
    x"FA",x"FD",x"5E",x"00",x"FD",x"56",x"01",x"FD", -- 0x1628
    x"6E",x"02",x"FD",x"66",x"03",x"F1",x"06",x"04", -- 0x1630
    x"CB",x"23",x"CB",x"12",x"ED",x"6A",x"10",x"F8", -- 0x1638
    x"FD",x"21",x"00",x"00",x"FD",x"39",x"FD",x"73", -- 0x1640
    x"00",x"FD",x"72",x"01",x"FD",x"75",x"02",x"FD", -- 0x1648
    x"74",x"03",x"21",x"16",x"00",x"39",x"EB",x"21", -- 0x1650
    x"0E",x"00",x"39",x"01",x"04",x"00",x"ED",x"B0", -- 0x1658
    x"AF",x"FD",x"21",x"04",x"00",x"FD",x"39",x"FD", -- 0x1660
    x"77",x"00",x"FD",x"77",x"01",x"FD",x"77",x"02", -- 0x1668
    x"FD",x"77",x"03",x"21",x"00",x"00",x"39",x"FD", -- 0x1670
    x"21",x"04",x"00",x"FD",x"39",x"FD",x"7E",x"00", -- 0x1678
    x"96",x"FD",x"7E",x"01",x"23",x"9E",x"FD",x"7E", -- 0x1680
    x"02",x"23",x"9E",x"FD",x"7E",x"03",x"23",x"9E", -- 0x1688
    x"D2",x"6B",x"18",x"FD",x"7E",x"00",x"E6",x"0F", -- 0x1690
    x"20",x"3B",x"FD",x"21",x"16",x"00",x"FD",x"39", -- 0x1698
    x"FD",x"4E",x"00",x"FD",x"46",x"01",x"FD",x"5E", -- 0x16A0
    x"02",x"FD",x"56",x"03",x"FD",x"34",x"00",x"20", -- 0x16A8
    x"0D",x"FD",x"34",x"01",x"20",x"08",x"FD",x"34", -- 0x16B0
    x"02",x"20",x"03",x"FD",x"34",x"03",x"21",x"55", -- 0x16B8
    x"FA",x"E5",x"D5",x"C5",x"CD",x"E8",x"07",x"F1", -- 0x16C0
    x"F1",x"F1",x"21",x"0C",x"00",x"39",x"36",x"55", -- 0x16C8
    x"23",x"36",x"FA",x"18",x"0D",x"21",x"0C",x"00", -- 0x16D0
    x"39",x"7E",x"C6",x"20",x"77",x"23",x"7E",x"CE", -- 0x16D8
    x"00",x"77",x"FD",x"21",x"0C",x"00",x"FD",x"39", -- 0x16E0
    x"FD",x"6E",x"00",x"FD",x"66",x"01",x"7E",x"B7", -- 0x16E8
    x"CA",x"4D",x"18",x"D6",x"E5",x"CA",x"4D",x"18", -- 0x16F0
    x"FD",x"6E",x"00",x"FD",x"66",x"01",x"11",x"0B", -- 0x16F8
    x"00",x"19",x"7E",x"E6",x"18",x"C2",x"4D",x"18", -- 0x1700
    x"21",x"0B",x"00",x"E5",x"21",x"26",x"00",x"39", -- 0x1708
    x"4E",x"23",x"46",x"C5",x"21",x"10",x"00",x"39", -- 0x1710
    x"4E",x"23",x"46",x"C5",x"CD",x"E2",x"0C",x"F1", -- 0x1718
    x"F1",x"F1",x"7C",x"B5",x"C2",x"4D",x"18",x"21", -- 0x1720
    x"22",x"00",x"39",x"7E",x"FD",x"21",x"14",x"00", -- 0x1728
    x"FD",x"39",x"FD",x"77",x"00",x"21",x"23",x"00", -- 0x1730
    x"39",x"7E",x"FD",x"21",x"14",x"00",x"FD",x"39", -- 0x1738
    x"FD",x"77",x"01",x"21",x"1E",x"00",x"39",x"FD", -- 0x1740
    x"7E",x"00",x"C6",x"04",x"77",x"FD",x"7E",x"01", -- 0x1748
    x"CE",x"00",x"23",x"77",x"21",x"0C",x"00",x"39", -- 0x1750
    x"7E",x"23",x"66",x"6F",x"11",x"1C",x"00",x"19", -- 0x1758
    x"4E",x"23",x"46",x"23",x"5E",x"23",x"56",x"21", -- 0x1760
    x"1E",x"00",x"39",x"7E",x"23",x"66",x"6F",x"71", -- 0x1768
    x"23",x"70",x"23",x"73",x"23",x"72",x"21",x"1E", -- 0x1770
    x"00",x"39",x"FD",x"21",x"14",x"00",x"FD",x"39", -- 0x1778
    x"FD",x"7E",x"00",x"C6",x"08",x"77",x"FD",x"7E", -- 0x1780
    x"01",x"CE",x"00",x"23",x"77",x"FD",x"21",x"0C", -- 0x1788
    x"00",x"FD",x"39",x"FD",x"6E",x"00",x"FD",x"66", -- 0x1790
    x"01",x"11",x"1A",x"00",x"19",x"7E",x"FD",x"21", -- 0x1798
    x"12",x"00",x"FD",x"39",x"FD",x"77",x"00",x"23", -- 0x17A0
    x"7E",x"FD",x"77",x"01",x"FD",x"21",x"2D",x"FA", -- 0x17A8
    x"FD",x"7E",x"01",x"FD",x"B6",x"00",x"28",x"40", -- 0x17B0
    x"21",x"0C",x"00",x"39",x"7E",x"23",x"66",x"6F", -- 0x17B8
    x"11",x"14",x"00",x"19",x"4E",x"23",x"7E",x"E6", -- 0x17C0
    x"0F",x"47",x"11",x"00",x"00",x"F5",x"FD",x"21", -- 0x17C8
    x"1C",x"00",x"FD",x"39",x"FD",x"71",x"00",x"FD", -- 0x17D0
    x"70",x"01",x"FD",x"73",x"02",x"FD",x"72",x"03", -- 0x17D8
    x"F1",x"3E",x"10",x"FD",x"CB",x"00",x"26",x"FD", -- 0x17E0
    x"CB",x"01",x"16",x"FD",x"CB",x"02",x"16",x"FD", -- 0x17E8
    x"CB",x"03",x"16",x"3D",x"20",x"ED",x"18",x"13", -- 0x17F0
    x"AF",x"FD",x"21",x"1A",x"00",x"FD",x"39",x"FD", -- 0x17F8
    x"77",x"00",x"FD",x"77",x"01",x"FD",x"77",x"02", -- 0x1800
    x"FD",x"77",x"03",x"21",x"12",x"00",x"39",x"4E", -- 0x1808
    x"23",x"46",x"11",x"00",x"00",x"79",x"21",x"1A", -- 0x1810
    x"00",x"39",x"86",x"4F",x"78",x"23",x"8E",x"47", -- 0x1818
    x"7B",x"23",x"8E",x"5F",x"7A",x"23",x"8E",x"57", -- 0x1820
    x"21",x"1E",x"00",x"39",x"7E",x"23",x"66",x"6F", -- 0x1828
    x"71",x"23",x"70",x"23",x"73",x"23",x"72",x"21", -- 0x1830
    x"14",x"00",x"39",x"7E",x"23",x"66",x"6F",x"AF", -- 0x1838
    x"77",x"23",x"77",x"23",x"AF",x"77",x"23",x"77", -- 0x1840
    x"2E",x"01",x"C3",x"67",x"19",x"FD",x"21",x"04", -- 0x1848
    x"00",x"FD",x"39",x"FD",x"34",x"00",x"C2",x"73", -- 0x1850
    x"16",x"FD",x"34",x"01",x"C2",x"73",x"16",x"FD", -- 0x1858
    x"34",x"02",x"C2",x"73",x"16",x"FD",x"34",x"03", -- 0x1860
    x"C3",x"73",x"16",x"FD",x"21",x"2D",x"FA",x"FD", -- 0x1868
    x"7E",x"01",x"FD",x"B6",x"00",x"CA",x"65",x"19", -- 0x1870
    x"FD",x"21",x"08",x"00",x"FD",x"39",x"FD",x"6E", -- 0x1878
    x"02",x"FD",x"66",x"03",x"E5",x"FD",x"6E",x"00", -- 0x1880
    x"FD",x"66",x"01",x"E5",x"CD",x"3A",x"0B",x"F1", -- 0x1888
    x"F1",x"FD",x"21",x"1A",x"00",x"FD",x"39",x"FD", -- 0x1890
    x"72",x"03",x"FD",x"73",x"02",x"FD",x"74",x"01", -- 0x1898
    x"FD",x"75",x"00",x"21",x"08",x"00",x"39",x"EB", -- 0x18A0
    x"21",x"1A",x"00",x"39",x"01",x"04",x"00",x"ED", -- 0x18A8
    x"B0",x"21",x"08",x"00",x"39",x"7E",x"E6",x"F8", -- 0x18B0
    x"FD",x"21",x"1A",x"00",x"FD",x"39",x"FD",x"77", -- 0x18B8
    x"00",x"21",x"09",x"00",x"39",x"7E",x"FD",x"21", -- 0x18C0
    x"1A",x"00",x"FD",x"39",x"FD",x"77",x"01",x"21", -- 0x18C8
    x"0A",x"00",x"39",x"7E",x"FD",x"21",x"1A",x"00", -- 0x18D0
    x"FD",x"39",x"FD",x"77",x"02",x"21",x"0B",x"00", -- 0x18D8
    x"39",x"7E",x"E6",x"0F",x"FD",x"21",x"1A",x"00", -- 0x18E0
    x"FD",x"39",x"FD",x"77",x"03",x"FD",x"7E",x"00", -- 0x18E8
    x"D6",x"F8",x"20",x"13",x"FD",x"7E",x"01",x"3C", -- 0x18F0
    x"20",x"0D",x"FD",x"7E",x"02",x"3C",x"20",x"07", -- 0x18F8
    x"FD",x"7E",x"03",x"D6",x"0F",x"28",x"5E",x"FD", -- 0x1900
    x"21",x"08",x"00",x"FD",x"39",x"FD",x"7E",x"00", -- 0x1908
    x"C6",x"FE",x"4F",x"FD",x"7E",x"01",x"CE",x"FF", -- 0x1910
    x"47",x"FD",x"7E",x"02",x"CE",x"FF",x"5F",x"FD", -- 0x1918
    x"7E",x"03",x"CE",x"FF",x"57",x"D5",x"C5",x"2A", -- 0x1920
    x"47",x"FA",x"E5",x"2A",x"45",x"FA",x"E5",x"CD", -- 0x1928
    x"7B",x"20",x"F1",x"F1",x"F1",x"F1",x"4D",x"44", -- 0x1930
    x"FD",x"21",x"33",x"FA",x"FD",x"7E",x"00",x"81", -- 0x1938
    x"4F",x"FD",x"7E",x"01",x"88",x"47",x"FD",x"7E", -- 0x1940
    x"02",x"8B",x"5F",x"FD",x"7E",x"03",x"8A",x"57", -- 0x1948
    x"FD",x"21",x"0E",x"00",x"FD",x"39",x"FD",x"71", -- 0x1950
    x"00",x"FD",x"70",x"01",x"FD",x"73",x"02",x"FD", -- 0x1958
    x"72",x"03",x"C3",x"52",x"16",x"2E",x"00",x"FD", -- 0x1960
    x"21",x"20",x"00",x"FD",x"39",x"FD",x"F9",x"C9", -- 0x1968
    x"21",x"F4",x"FF",x"39",x"F9",x"21",x"08",x"00", -- 0x1970
    x"39",x"EB",x"21",x"33",x"FA",x"01",x"04",x"00", -- 0x1978
    x"ED",x"B0",x"21",x"0E",x"00",x"39",x"7E",x"FD", -- 0x1980
    x"21",x"06",x"00",x"FD",x"39",x"FD",x"77",x"00", -- 0x1988
    x"21",x"0F",x"00",x"39",x"7E",x"FD",x"21",x"06", -- 0x1990
    x"00",x"FD",x"39",x"FD",x"77",x"01",x"21",x"04", -- 0x1998
    x"00",x"39",x"FD",x"7E",x"00",x"C6",x"08",x"77", -- 0x19A0
    x"FD",x"7E",x"01",x"CE",x"00",x"23",x"77",x"21", -- 0x19A8
    x"04",x"00",x"39",x"7E",x"23",x"66",x"6F",x"4E", -- 0x19B0
    x"23",x"46",x"23",x"5E",x"23",x"56",x"79",x"C6", -- 0x19B8
    x"FE",x"4F",x"78",x"CE",x"FF",x"47",x"7B",x"CE", -- 0x19C0
    x"FF",x"5F",x"7A",x"CE",x"FF",x"57",x"D5",x"C5", -- 0x19C8
    x"2A",x"47",x"FA",x"E5",x"2A",x"45",x"FA",x"E5", -- 0x19D0
    x"CD",x"7B",x"20",x"F1",x"F1",x"F1",x"F1",x"4D", -- 0x19D8
    x"44",x"FD",x"21",x"08",x"00",x"FD",x"39",x"FD", -- 0x19E0
    x"7E",x"00",x"81",x"4F",x"FD",x"7E",x"01",x"88", -- 0x19E8
    x"47",x"FD",x"7E",x"02",x"8B",x"5F",x"FD",x"7E", -- 0x19F0
    x"03",x"8A",x"57",x"FD",x"21",x"00",x"00",x"FD", -- 0x19F8
    x"39",x"FD",x"71",x"00",x"FD",x"70",x"01",x"FD", -- 0x1A00
    x"73",x"02",x"FD",x"72",x"03",x"21",x"06",x"00", -- 0x1A08
    x"39",x"7E",x"23",x"66",x"6F",x"4E",x"23",x"46", -- 0x1A10
    x"23",x"5E",x"23",x"56",x"79",x"FD",x"21",x"49", -- 0x1A18
    x"FA",x"FD",x"A6",x"00",x"4F",x"78",x"FD",x"A6", -- 0x1A20
    x"01",x"47",x"7B",x"FD",x"A6",x"02",x"5F",x"7A", -- 0x1A28
    x"FD",x"A6",x"03",x"57",x"FD",x"21",x"00",x"00", -- 0x1A30
    x"FD",x"39",x"FD",x"7E",x"00",x"81",x"4F",x"FD", -- 0x1A38
    x"7E",x"01",x"88",x"47",x"FD",x"7E",x"02",x"8B", -- 0x1A40
    x"5F",x"FD",x"7E",x"03",x"8A",x"57",x"21",x"10", -- 0x1A48
    x"00",x"39",x"7E",x"23",x"66",x"6F",x"E5",x"D5", -- 0x1A50
    x"C5",x"CD",x"E8",x"07",x"F1",x"F1",x"F1",x"7D", -- 0x1A58
    x"B7",x"20",x"03",x"6F",x"18",x"6F",x"FD",x"21", -- 0x1A60
    x"06",x"00",x"FD",x"39",x"FD",x"6E",x"00",x"FD", -- 0x1A68
    x"66",x"01",x"4E",x"23",x"46",x"23",x"5E",x"23", -- 0x1A70
    x"56",x"0C",x"20",x"07",x"04",x"20",x"04",x"1C", -- 0x1A78
    x"20",x"01",x"14",x"FD",x"6E",x"00",x"FD",x"66", -- 0x1A80
    x"01",x"71",x"23",x"70",x"23",x"73",x"23",x"72", -- 0x1A88
    x"79",x"FD",x"21",x"49",x"FA",x"FD",x"A6",x"00", -- 0x1A90
    x"4F",x"78",x"FD",x"A6",x"01",x"47",x"7B",x"FD", -- 0x1A98
    x"A6",x"02",x"5F",x"7A",x"FD",x"A6",x"03",x"B3", -- 0x1AA0
    x"B0",x"B1",x"20",x"27",x"21",x"04",x"00",x"39", -- 0x1AA8
    x"7E",x"23",x"66",x"6F",x"4E",x"23",x"46",x"23", -- 0x1AB0
    x"5E",x"23",x"56",x"D5",x"C5",x"CD",x"3A",x"0B", -- 0x1AB8
    x"F1",x"F1",x"4D",x"44",x"21",x"04",x"00",x"39", -- 0x1AC0
    x"7E",x"23",x"66",x"6F",x"71",x"23",x"70",x"23", -- 0x1AC8
    x"73",x"23",x"72",x"2E",x"01",x"FD",x"21",x"0C", -- 0x1AD0
    x"00",x"FD",x"39",x"FD",x"F9",x"C9",x"3E",x"40", -- 0x1AD8
    x"01",x"3B",x"24",x"ED",x"79",x"3E",x"00",x"01", -- 0x1AE0
    x"3B",x"25",x"ED",x"79",x"3E",x"41",x"01",x"3B", -- 0x1AE8
    x"24",x"ED",x"79",x"01",x"00",x"00",x"C5",x"79", -- 0x1AF0
    x"01",x"3B",x"25",x"ED",x"79",x"C1",x"03",x"78", -- 0x1AF8
    x"D6",x"01",x"38",x"F2",x"C9",x"00",x"00",x"00", -- 0x1B00
    x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10", -- 0x1B08
    x"10",x"10",x"00",x"10",x"00",x"00",x"24",x"24", -- 0x1B10
    x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"7E", -- 0x1B18
    x"24",x"24",x"7E",x"24",x"00",x"00",x"08",x"3E", -- 0x1B20
    x"28",x"3E",x"0A",x"3E",x"08",x"00",x"62",x"64", -- 0x1B28
    x"08",x"10",x"26",x"46",x"00",x"00",x"10",x"28", -- 0x1B30
    x"10",x"2A",x"44",x"3A",x"00",x"00",x"08",x"10", -- 0x1B38
    x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08", -- 0x1B40
    x"08",x"08",x"08",x"04",x"00",x"00",x"20",x"10", -- 0x1B48
    x"10",x"10",x"10",x"20",x"00",x"00",x"00",x"14", -- 0x1B50
    x"08",x"3E",x"08",x"14",x"00",x"00",x"00",x"08", -- 0x1B58
    x"08",x"3E",x"08",x"08",x"00",x"00",x"00",x"00", -- 0x1B60
    x"00",x"00",x"08",x"08",x"10",x"00",x"00",x"00", -- 0x1B68
    x"00",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B70
    x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"02", -- 0x1B78
    x"04",x"08",x"10",x"20",x"00",x"00",x"3C",x"46", -- 0x1B80
    x"4A",x"52",x"62",x"3C",x"00",x"00",x"18",x"28", -- 0x1B88
    x"08",x"08",x"08",x"3E",x"00",x"00",x"3C",x"42", -- 0x1B90
    x"02",x"3C",x"40",x"7E",x"00",x"00",x"3C",x"42", -- 0x1B98
    x"0C",x"02",x"42",x"3C",x"00",x"00",x"08",x"18", -- 0x1BA0
    x"28",x"48",x"7E",x"08",x"00",x"00",x"7E",x"40", -- 0x1BA8
    x"7C",x"02",x"42",x"3C",x"00",x"00",x"3C",x"40", -- 0x1BB0
    x"7C",x"42",x"42",x"3C",x"00",x"00",x"7E",x"02", -- 0x1BB8
    x"04",x"08",x"10",x"10",x"00",x"00",x"3C",x"42", -- 0x1BC0
    x"3C",x"42",x"42",x"3C",x"00",x"00",x"3C",x"42", -- 0x1BC8
    x"42",x"3E",x"02",x"3C",x"00",x"00",x"00",x"00", -- 0x1BD0
    x"10",x"00",x"00",x"10",x"00",x"00",x"00",x"10", -- 0x1BD8
    x"00",x"00",x"10",x"10",x"20",x"00",x"00",x"04", -- 0x1BE0
    x"08",x"10",x"08",x"04",x"00",x"00",x"00",x"00", -- 0x1BE8
    x"3E",x"00",x"3E",x"00",x"00",x"00",x"00",x"20", -- 0x1BF0
    x"10",x"08",x"10",x"20",x"00",x"00",x"3C",x"42", -- 0x1BF8
    x"04",x"08",x"00",x"08",x"00",x"00",x"3C",x"4A", -- 0x1C00
    x"56",x"5E",x"40",x"3C",x"00",x"00",x"3C",x"42", -- 0x1C08
    x"42",x"7E",x"42",x"42",x"00",x"00",x"7C",x"42", -- 0x1C10
    x"7C",x"42",x"42",x"7C",x"00",x"00",x"3C",x"42", -- 0x1C18
    x"40",x"40",x"42",x"3C",x"00",x"00",x"78",x"44", -- 0x1C20
    x"42",x"42",x"44",x"78",x"00",x"00",x"7E",x"40", -- 0x1C28
    x"7C",x"40",x"40",x"7E",x"00",x"00",x"7E",x"40", -- 0x1C30
    x"7C",x"40",x"40",x"40",x"00",x"00",x"3C",x"42", -- 0x1C38
    x"40",x"4E",x"42",x"3C",x"00",x"00",x"42",x"42", -- 0x1C40
    x"7E",x"42",x"42",x"42",x"00",x"00",x"3E",x"08", -- 0x1C48
    x"08",x"08",x"08",x"3E",x"00",x"00",x"02",x"02", -- 0x1C50
    x"02",x"42",x"42",x"3C",x"00",x"00",x"44",x"48", -- 0x1C58
    x"70",x"48",x"44",x"42",x"00",x"00",x"40",x"40", -- 0x1C60
    x"40",x"40",x"40",x"7E",x"00",x"00",x"42",x"66", -- 0x1C68
    x"5A",x"42",x"42",x"42",x"00",x"00",x"42",x"62", -- 0x1C70
    x"52",x"4A",x"46",x"42",x"00",x"00",x"3C",x"42", -- 0x1C78
    x"42",x"42",x"42",x"3C",x"00",x"00",x"7C",x"42", -- 0x1C80
    x"42",x"7C",x"40",x"40",x"00",x"00",x"3C",x"42", -- 0x1C88
    x"42",x"52",x"4A",x"3C",x"00",x"00",x"7C",x"42", -- 0x1C90
    x"42",x"7C",x"44",x"42",x"00",x"00",x"3C",x"40", -- 0x1C98
    x"3C",x"02",x"42",x"3C",x"00",x"00",x"FE",x"10", -- 0x1CA0
    x"10",x"10",x"10",x"10",x"00",x"00",x"42",x"42", -- 0x1CA8
    x"42",x"42",x"42",x"3C",x"00",x"00",x"42",x"42", -- 0x1CB0
    x"42",x"42",x"24",x"18",x"00",x"00",x"42",x"42", -- 0x1CB8
    x"42",x"42",x"5A",x"24",x"00",x"00",x"42",x"24", -- 0x1CC0
    x"18",x"18",x"24",x"42",x"00",x"00",x"82",x"44", -- 0x1CC8
    x"28",x"10",x"10",x"10",x"00",x"00",x"7E",x"04", -- 0x1CD0
    x"08",x"10",x"20",x"7E",x"00",x"00",x"0E",x"08", -- 0x1CD8
    x"08",x"08",x"08",x"0E",x"00",x"00",x"00",x"40", -- 0x1CE0
    x"20",x"10",x"08",x"04",x"00",x"00",x"70",x"10", -- 0x1CE8
    x"10",x"10",x"10",x"70",x"00",x"00",x"10",x"38", -- 0x1CF0
    x"54",x"10",x"10",x"10",x"00",x"00",x"00",x"00", -- 0x1CF8
    x"00",x"00",x"00",x"00",x"FF",x"00",x"1C",x"22", -- 0x1D00
    x"78",x"20",x"20",x"7E",x"00",x"00",x"00",x"38", -- 0x1D08
    x"04",x"3C",x"44",x"3C",x"00",x"00",x"20",x"20", -- 0x1D10
    x"3C",x"22",x"22",x"3C",x"00",x"00",x"00",x"1C", -- 0x1D18
    x"20",x"20",x"20",x"1C",x"00",x"00",x"04",x"04", -- 0x1D20
    x"3C",x"44",x"44",x"3C",x"00",x"00",x"00",x"38", -- 0x1D28
    x"44",x"78",x"40",x"3C",x"00",x"00",x"0C",x"10", -- 0x1D30
    x"18",x"10",x"10",x"10",x"00",x"00",x"00",x"3C", -- 0x1D38
    x"44",x"44",x"3C",x"04",x"38",x"00",x"40",x"40", -- 0x1D40
    x"78",x"44",x"44",x"44",x"00",x"00",x"10",x"00", -- 0x1D48
    x"30",x"10",x"10",x"38",x"00",x"00",x"04",x"00", -- 0x1D50
    x"04",x"04",x"04",x"24",x"18",x"00",x"20",x"28", -- 0x1D58
    x"30",x"30",x"28",x"24",x"00",x"00",x"10",x"10", -- 0x1D60
    x"10",x"10",x"10",x"0C",x"00",x"00",x"00",x"68", -- 0x1D68
    x"54",x"54",x"54",x"54",x"00",x"00",x"00",x"78", -- 0x1D70
    x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"38", -- 0x1D78
    x"44",x"44",x"44",x"38",x"00",x"00",x"00",x"78", -- 0x1D80
    x"44",x"44",x"78",x"40",x"40",x"00",x"00",x"3C", -- 0x1D88
    x"44",x"44",x"3C",x"04",x"06",x"00",x"00",x"1C", -- 0x1D90
    x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"38", -- 0x1D98
    x"40",x"38",x"04",x"78",x"00",x"00",x"10",x"38", -- 0x1DA0
    x"10",x"10",x"10",x"0C",x"00",x"00",x"00",x"44", -- 0x1DA8
    x"44",x"44",x"44",x"38",x"00",x"00",x"00",x"44", -- 0x1DB0
    x"44",x"28",x"28",x"10",x"00",x"00",x"00",x"44", -- 0x1DB8
    x"54",x"54",x"54",x"28",x"00",x"00",x"00",x"44", -- 0x1DC0
    x"28",x"10",x"28",x"44",x"00",x"00",x"00",x"44", -- 0x1DC8
    x"44",x"44",x"3C",x"04",x"38",x"00",x"00",x"7C", -- 0x1DD0
    x"08",x"10",x"20",x"7C",x"00",x"00",x"0E",x"08", -- 0x1DD8
    x"30",x"08",x"08",x"0E",x"00",x"00",x"08",x"08", -- 0x1DE0
    x"08",x"08",x"08",x"08",x"00",x"00",x"70",x"10", -- 0x1DE8
    x"0C",x"10",x"10",x"70",x"00",x"00",x"14",x"28", -- 0x1DF0
    x"00",x"00",x"00",x"00",x"00",x"3C",x"42",x"99", -- 0x1DF8
    x"A1",x"A1",x"99",x"42",x"3C",x"21",x"62",x"FC", -- 0x1E00
    x"36",x"00",x"21",x"61",x"FC",x"36",x"00",x"01", -- 0x1E08
    x"00",x"40",x"59",x"50",x"AF",x"12",x"03",x"78", -- 0x1E10
    x"D6",x"58",x"38",x"F6",x"01",x"00",x"58",x"69", -- 0x1E18
    x"60",x"36",x"47",x"03",x"78",x"D6",x"5B",x"38", -- 0x1E20
    x"F6",x"C9",x"21",x"02",x"00",x"39",x"7E",x"E6", -- 0x1E28
    x"1F",x"32",x"61",x"FC",x"21",x"03",x"00",x"39", -- 0x1E30
    x"7E",x"FD",x"21",x"62",x"FC",x"FD",x"77",x"00", -- 0x1E38
    x"3E",x"17",x"FD",x"96",x"00",x"D0",x"FD",x"36", -- 0x1E40
    x"00",x"17",x"C9",x"F5",x"F5",x"21",x"06",x"00", -- 0x1E48
    x"39",x"7E",x"D6",x"0A",x"20",x"1B",x"21",x"61", -- 0x1E50
    x"FC",x"36",x"00",x"FD",x"21",x"62",x"FC",x"FD", -- 0x1E58
    x"34",x"00",x"3E",x"17",x"FD",x"96",x"00",x"D2", -- 0x1E60
    x"B1",x"1F",x"FD",x"36",x"00",x"17",x"C3",x"B1", -- 0x1E68
    x"1F",x"21",x"06",x"00",x"39",x"7E",x"D6",x"08", -- 0x1E70
    x"20",x"26",x"FD",x"21",x"61",x"FC",x"FD",x"7E", -- 0x1E78
    x"00",x"B7",x"20",x"15",x"FD",x"36",x"00",x"1F", -- 0x1E80
    x"FD",x"21",x"62",x"FC",x"FD",x"7E",x"00",x"B7", -- 0x1E88
    x"CA",x"B1",x"1F",x"FD",x"35",x"00",x"C3",x"B1", -- 0x1E90
    x"1F",x"21",x"61",x"FC",x"35",x"C3",x"B1",x"1F", -- 0x1E98
    x"21",x"06",x"00",x"39",x"7E",x"06",x"00",x"C6", -- 0x1EA0
    x"E0",x"4F",x"78",x"CE",x"FF",x"47",x"CB",x"21", -- 0x1EA8
    x"CB",x"10",x"CB",x"21",x"CB",x"10",x"CB",x"21", -- 0x1EB0
    x"CB",x"10",x"ED",x"43",x"5B",x"FC",x"3A",x"62", -- 0x1EB8
    x"FC",x"FD",x"21",x"00",x"00",x"FD",x"39",x"FD", -- 0x1EC0
    x"77",x"00",x"FD",x"36",x"01",x"00",x"FD",x"7E", -- 0x1EC8
    x"00",x"FD",x"21",x"5D",x"FC",x"FD",x"77",x"01", -- 0x1ED0
    x"FD",x"36",x"00",x"00",x"0E",x"00",x"FD",x"7E", -- 0x1ED8
    x"01",x"E6",x"18",x"47",x"FD",x"7E",x"00",x"E6", -- 0x1EE0
    x"E0",x"6F",x"26",x"00",x"29",x"29",x"29",x"79", -- 0x1EE8
    x"B5",x"4F",x"78",x"B4",x"47",x"1E",x"00",x"FD", -- 0x1EF0
    x"7E",x"01",x"E6",x"07",x"57",x"3E",x"03",x"CB", -- 0x1EF8
    x"3A",x"CB",x"1B",x"3D",x"20",x"F9",x"79",x"B3", -- 0x1F00
    x"FD",x"77",x"00",x"78",x"B2",x"FD",x"77",x"01", -- 0x1F08
    x"FD",x"7E",x"00",x"C6",x"00",x"5F",x"FD",x"7E", -- 0x1F10
    x"01",x"CE",x"40",x"57",x"21",x"61",x"FC",x"4E", -- 0x1F18
    x"06",x"00",x"FD",x"21",x"02",x"00",x"FD",x"39", -- 0x1F20
    x"FD",x"71",x"00",x"FD",x"70",x"01",x"7B",x"21", -- 0x1F28
    x"02",x"00",x"39",x"FD",x"21",x"5D",x"FC",x"86", -- 0x1F30
    x"FD",x"77",x"00",x"7A",x"23",x"8E",x"FD",x"23", -- 0x1F38
    x"FD",x"77",x"00",x"E1",x"E5",x"29",x"29",x"29", -- 0x1F40
    x"29",x"29",x"5D",x"7C",x"C6",x"58",x"57",x"7B", -- 0x1F48
    x"21",x"5F",x"FC",x"81",x"77",x"7A",x"88",x"23", -- 0x1F50
    x"77",x"0E",x"00",x"ED",x"5B",x"5D",x"FC",x"FD", -- 0x1F58
    x"21",x"05",x"1B",x"C5",x"ED",x"4B",x"5B",x"FC", -- 0x1F60
    x"FD",x"09",x"C1",x"FD",x"7E",x"00",x"12",x"21", -- 0x1F68
    x"5D",x"FC",x"7E",x"C6",x"00",x"77",x"23",x"7E", -- 0x1F70
    x"CE",x"01",x"77",x"FD",x"21",x"5B",x"FC",x"FD", -- 0x1F78
    x"34",x"00",x"20",x"03",x"FD",x"34",x"01",x"0C", -- 0x1F80
    x"79",x"D6",x"08",x"38",x"CE",x"FD",x"21",x"61", -- 0x1F88
    x"FC",x"FD",x"34",x"00",x"3E",x"1F",x"FD",x"96", -- 0x1F90
    x"00",x"30",x"16",x"FD",x"36",x"00",x"00",x"FD", -- 0x1F98
    x"21",x"62",x"FC",x"FD",x"34",x"00",x"3E",x"17", -- 0x1FA0
    x"FD",x"96",x"00",x"30",x"04",x"FD",x"36",x"00", -- 0x1FA8
    x"17",x"F1",x"F1",x"C9",x"D1",x"C1",x"C5",x"D5", -- 0x1FB0
    x"0A",x"03",x"57",x"B7",x"C8",x"C5",x"D5",x"33", -- 0x1FB8
    x"CD",x"4B",x"1E",x"33",x"C1",x"18",x"F1",x"21", -- 0x1FC0
    x"F0",x"FF",x"39",x"F9",x"21",x"00",x"00",x"39", -- 0x1FC8
    x"4D",x"44",x"36",x"30",x"69",x"60",x"23",x"36", -- 0x1FD0
    x"31",x"69",x"60",x"23",x"23",x"36",x"32",x"69", -- 0x1FD8
    x"60",x"23",x"23",x"23",x"36",x"33",x"21",x"04", -- 0x1FE0
    x"00",x"09",x"36",x"34",x"21",x"05",x"00",x"09", -- 0x1FE8
    x"36",x"35",x"21",x"06",x"00",x"09",x"36",x"36", -- 0x1FF0
    x"21",x"07",x"00",x"09",x"36",x"37",x"21",x"08", -- 0x1FF8
    x"00",x"09",x"36",x"38",x"21",x"09",x"00",x"09", -- 0x2000
    x"36",x"39",x"21",x"0A",x"00",x"09",x"36",x"41", -- 0x2008
    x"21",x"0B",x"00",x"09",x"36",x"42",x"21",x"0C", -- 0x2010
    x"00",x"09",x"36",x"43",x"21",x"0D",x"00",x"09", -- 0x2018
    x"36",x"44",x"21",x"0E",x"00",x"09",x"36",x"45", -- 0x2020
    x"21",x"0F",x"00",x"09",x"36",x"46",x"21",x"12", -- 0x2028
    x"00",x"39",x"7E",x"E6",x"F0",x"07",x"07",x"07", -- 0x2030
    x"07",x"E6",x"0F",x"5F",x"6B",x"26",x"00",x"09", -- 0x2038
    x"56",x"C5",x"D5",x"33",x"CD",x"4B",x"1E",x"33", -- 0x2040
    x"C1",x"21",x"12",x"00",x"39",x"7E",x"E6",x"0F", -- 0x2048
    x"6F",x"26",x"00",x"09",x"46",x"C5",x"33",x"CD", -- 0x2050
    x"4B",x"1E",x"33",x"21",x"10",x"00",x"39",x"F9", -- 0x2058
    x"C9",x"F1",x"C1",x"D1",x"D5",x"C5",x"F5",x"AF", -- 0x2060
    x"6F",x"B0",x"06",x"10",x"20",x"04",x"06",x"08", -- 0x2068
    x"79",x"29",x"CB",x"11",x"17",x"30",x"01",x"19", -- 0x2070
    x"10",x"F7",x"C9",x"DD",x"E5",x"DD",x"21",x"00", -- 0x2078
    x"00",x"DD",x"39",x"21",x"FA",x"FF",x"39",x"F9", -- 0x2080
    x"21",x"0A",x"00",x"39",x"EB",x"4B",x"42",x"03", -- 0x2088
    x"03",x"DD",x"71",x"FE",x"DD",x"70",x"FF",x"6B", -- 0x2090
    x"62",x"23",x"23",x"4E",x"23",x"46",x"21",x"0E", -- 0x2098
    x"00",x"39",x"DD",x"75",x"FC",x"DD",x"74",x"FD", -- 0x20A0
    x"DD",x"6E",x"FC",x"DD",x"66",x"FD",x"7E",x"23", -- 0x20A8
    x"66",x"6F",x"D5",x"E5",x"C5",x"CD",x"61",x"20", -- 0x20B0
    x"F1",x"F1",x"4D",x"44",x"D1",x"DD",x"6E",x"FE", -- 0x20B8
    x"DD",x"66",x"FF",x"71",x"23",x"70",x"4B",x"42", -- 0x20C0
    x"03",x"03",x"DD",x"71",x"FE",x"DD",x"70",x"FF", -- 0x20C8
    x"6B",x"62",x"23",x"23",x"7E",x"DD",x"77",x"FA", -- 0x20D0
    x"23",x"7E",x"DD",x"77",x"FB",x"C1",x"E1",x"E5", -- 0x20D8
    x"C5",x"23",x"23",x"4E",x"23",x"46",x"6B",x"62", -- 0x20E0
    x"7E",x"23",x"66",x"6F",x"D5",x"E5",x"C5",x"CD", -- 0x20E8
    x"61",x"20",x"F1",x"F1",x"D1",x"DD",x"7E",x"FA", -- 0x20F0
    x"85",x"4F",x"DD",x"7E",x"FB",x"8C",x"47",x"DD", -- 0x20F8
    x"6E",x"FE",x"DD",x"66",x"FF",x"71",x"23",x"70", -- 0x2100
    x"4B",x"42",x"03",x"03",x"33",x"33",x"C5",x"6B", -- 0x2108
    x"62",x"23",x"23",x"4E",x"23",x"46",x"6B",x"62", -- 0x2110
    x"23",x"7E",x"DD",x"77",x"FE",x"DD",x"6E",x"FC", -- 0x2118
    x"DD",x"66",x"FD",x"23",x"66",x"D5",x"C5",x"DD", -- 0x2120
    x"5E",x"FE",x"2E",x"00",x"55",x"06",x"08",x"29", -- 0x2128
    x"30",x"01",x"19",x"10",x"FA",x"C1",x"D1",x"09", -- 0x2130
    x"4D",x"44",x"E1",x"E5",x"71",x"23",x"70",x"C1", -- 0x2138
    x"E1",x"E5",x"C5",x"4E",x"6B",x"62",x"23",x"66", -- 0x2140
    x"D5",x"59",x"2E",x"00",x"55",x"06",x"08",x"29", -- 0x2148
    x"30",x"01",x"19",x"10",x"FA",x"D1",x"4D",x"44", -- 0x2150
    x"DD",x"6E",x"FC",x"DD",x"66",x"FD",x"23",x"E5", -- 0x2158
    x"FD",x"E1",x"6B",x"62",x"7E",x"DD",x"77",x"FA", -- 0x2160
    x"DD",x"6E",x"FC",x"DD",x"66",x"FD",x"23",x"6E", -- 0x2168
    x"D5",x"C5",x"5D",x"DD",x"66",x"FA",x"2E",x"00", -- 0x2170
    x"55",x"06",x"08",x"29",x"30",x"01",x"19",x"10", -- 0x2178
    x"FA",x"C1",x"D1",x"FD",x"75",x"00",x"FD",x"74", -- 0x2180
    x"01",x"DD",x"6E",x"FC",x"DD",x"66",x"FD",x"23", -- 0x2188
    x"23",x"23",x"E3",x"DD",x"6E",x"FC",x"DD",x"66", -- 0x2190
    x"FD",x"23",x"E5",x"FD",x"E1",x"DD",x"6E",x"FC", -- 0x2198
    x"DD",x"66",x"FD",x"23",x"7E",x"23",x"66",x"6F", -- 0x21A0
    x"09",x"FD",x"75",x"00",x"FD",x"74",x"01",x"BF", -- 0x21A8
    x"ED",x"42",x"3E",x"00",x"17",x"E1",x"E5",x"77", -- 0x21B0
    x"4B",x"42",x"1A",x"5F",x"DD",x"6E",x"FC",x"DD", -- 0x21B8
    x"66",x"FD",x"66",x"C5",x"2E",x"00",x"55",x"06", -- 0x21C0
    x"08",x"29",x"30",x"01",x"19",x"10",x"FA",x"C1", -- 0x21C8
    x"EB",x"7B",x"02",x"03",x"7A",x"02",x"D1",x"C1", -- 0x21D0
    x"C5",x"D5",x"AF",x"02",x"DD",x"7E",x"04",x"DD", -- 0x21D8
    x"86",x"08",x"6F",x"DD",x"7E",x"05",x"DD",x"8E", -- 0x21E0
    x"09",x"67",x"DD",x"7E",x"06",x"DD",x"8E",x"0A", -- 0x21E8
    x"5F",x"DD",x"7E",x"07",x"DD",x"8E",x"0B",x"57", -- 0x21F0
    x"DD",x"F9",x"DD",x"E1",x"C9",x"5E",x"07",x"00", -- 0x21F8
    x"01",x"03",x"00",x"78",x"B1",x"28",x"08",x"11", -- 0x2200
    x"63",x"FC",x"21",x"FD",x"21",x"ED",x"B0",x"C9", -- 0x2208
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2210
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2218
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2220
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2228
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2230
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2238
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2240
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2248
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2250
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2258
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2260
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2268
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2270
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2278
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2280
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2288
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2290
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2298
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2300
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2308
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2310
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2318
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2320
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2328
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2330
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2338
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2340
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2348
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2350
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2358
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2360
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2368
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2370
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2378
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2380
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2388
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2390
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2398
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2400
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2408
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2410
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2418
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2420
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2428
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2430
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2438
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2440
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2448
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2450
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2458
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2460
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2468
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2470
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2478
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2480
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2488
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2490
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2498
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2500
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2508
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2510
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2518
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2520
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2528
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2530
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2538
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2540
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2548
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2550
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2558
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2560
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2568
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2570
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2578
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2580
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2588
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2590
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2598
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2600
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2608
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2610
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2618
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2620
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2628
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2630
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2638
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2640
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2648
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2650
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2658
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2660
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2668
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2670
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2678
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2680
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2688
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2690
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2698
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2700
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2708
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2710
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2718
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2720
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2728
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2730
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2738
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2740
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2748
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2750
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2758
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2760
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2768
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2770
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2778
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2780
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2788
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2790
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2798
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2800
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2808
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2810
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2818
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2820
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2828
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2830
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2838
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2840
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2848
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2850
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2858
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2860
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2868
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2870
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2878
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2880
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2888
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2890
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2898
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2900
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2908
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2910
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2918
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2920
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2928
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2930
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2938
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2940
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2948
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2950
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2958
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2960
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2968
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2970
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2978
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2980
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2988
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2990
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2998
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2ED0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2ED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3000
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3008
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3010
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3018
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3020
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3028
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3030
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3038
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3040
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3048
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3050
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3060
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3068
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3070
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3078
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3080
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3088
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3090
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3098
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3100
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3108
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3110
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3118
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3120
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3128
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3130
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3138
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3140
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3148
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3150
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3158
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3160
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3168
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3170
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3178
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3180
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3188
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3190
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3198
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3200
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3208
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3210
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3218
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3220
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3228
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3230
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3238
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3240
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3248
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3250
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3258
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3260
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3268
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3270
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3278
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3280
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3288
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3290
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3298
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3300
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3308
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3310
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3318
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3320
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3328
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3330
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3338
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3340
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3348
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3350
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3358
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3360
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3368
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3370
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3378
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3380
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3388
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3390
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3398
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3400
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3408
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3410
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3418
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3420
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3428
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3430
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3438
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3440
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3448
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3450
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3458
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3460
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3468
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3470
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3478
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3480
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3488
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3490
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3498
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3500
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3508
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3510
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3518
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3520
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3528
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3530
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3538
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3540
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3548
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3550
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3558
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3560
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3568
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3570
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3578
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3580
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3588
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3590
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3598
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3600
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3608
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3610
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3618
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3620
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3628
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3630
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3638
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3640
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3648
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3650
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3658
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3660
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3668
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3670
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3678
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3680
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3688
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3690
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3698
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3700
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3708
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3710
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3718
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3720
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3728
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3730
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3738
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3740
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3748
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3750
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3758
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3760
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3768
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3770
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3778
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3780
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3788
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3790
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3798
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3800
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3808
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3810
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3818
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3820
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3828
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3830
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3838
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3840
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3848
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3850
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3858
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3860
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3868
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3870
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3878
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3880
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3888
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3890
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3898
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3900
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3908
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3910
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3918
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3920
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3928
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3930
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3938
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3940
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3948
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3950
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3958
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3960
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3968
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3970
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3978
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3980
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3988
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3990
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3998
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x39F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3ED0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3ED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x3FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
